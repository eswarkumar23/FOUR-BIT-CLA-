magic
tech scmos
timestamp 1731666753
<< nwell >>
rect 0 0 34 24
rect 40 -1 64 23
<< ntransistor >>
rect 11 -26 13 -14
rect 21 -26 23 -14
rect 51 -15 53 -9
<< ptransistor >>
rect 11 6 13 18
rect 21 6 23 18
rect 51 5 53 17
<< ndiffusion >>
rect 10 -26 11 -14
rect 13 -26 21 -14
rect 23 -26 24 -14
rect 50 -15 51 -9
rect 53 -15 54 -9
<< pdiffusion >>
rect 10 6 11 18
rect 13 6 15 18
rect 19 6 21 18
rect 23 6 24 18
rect 50 5 51 17
rect 53 5 54 17
<< ndcontact >>
rect 6 -26 10 -14
rect 24 -26 28 -14
rect 46 -15 50 -9
rect 54 -15 58 -9
<< pdcontact >>
rect 6 6 10 18
rect 15 6 19 18
rect 24 6 28 18
rect 46 5 50 17
rect 54 5 58 17
<< polysilicon >>
rect 11 18 13 21
rect 21 18 23 21
rect 51 17 53 20
rect 11 -14 13 6
rect 21 -14 23 6
rect 51 -9 53 5
rect 51 -18 53 -15
rect 11 -29 13 -26
rect 21 -29 23 -26
<< polycontact >>
rect 7 -5 11 -1
rect 17 -11 21 -7
rect 47 -6 51 -2
<< metal1 >>
rect 0 26 43 27
rect 0 24 64 26
rect 6 18 9 24
rect 25 18 28 24
rect 40 23 64 24
rect 46 17 49 23
rect 15 3 18 6
rect 15 0 28 3
rect 0 -5 7 -2
rect 25 -3 28 0
rect 25 -6 47 -3
rect 55 -3 58 5
rect 55 -6 64 -3
rect 0 -11 17 -8
rect 25 -14 28 -6
rect 55 -9 58 -6
rect 46 -19 49 -15
rect 36 -22 64 -19
rect 6 -32 9 -26
rect 36 -32 40 -22
rect 0 -35 40 -32
<< labels >>
rlabel metal1 24 26 24 26 5 vdd!
rlabel metal1 24 -34 24 -34 1 gnd!
rlabel metal1 0 -11 0 -8 3 b
rlabel metal1 34 -6 34 -3 7 out
rlabel metal1 0 -5 0 -2 3 a
rlabel metal1 54 24 54 24 5 vdd!
rlabel metal1 60 -21 60 -21 1 gnd!
rlabel metal1 40 -6 40 -3 3 in
rlabel metal1 64 -6 64 -3 7 op
<< end >>
