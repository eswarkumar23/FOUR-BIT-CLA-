.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd
.option scale=0.09u
Vdd    vdd gnd 'SUPPLY'
vin    A 0 pulse 0 1.8 0ns 0ns 0ns 10ns 20ns
vin2   B 0 pulse 0 1.8 0ns 0ns 0ns 22ns 44ns 

M1000 a_n85_n22# A GND Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=200 ps=100
M1001 a_n85_n22# A VDD w_n98_8# CMOSP w=40 l=2
+  ad=200 pd=90 as=400 ps=180
M1002 B A out w_n28_13# CMOSP w=20 l=2
+  ad=100 pd=50 as=200 ps=100
M1003 a_n55_n10# B VDD w_15_7# CMOSP w=40 l=2
+  ad=300 pd=140 as=0 ps=0
M1004 a_n55_n10# B GND Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1005 out a_n85_n22# a_n55_n10# w_n61_n20# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 out A a_n55_n10# Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1007 B a_n85_n22# out Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 a_n55_n10# w_n61_n20# 0.06fF
C1 a_n55_n10# VDD 0.51fF
C2 a_n85_n22# A 0.07fF
C3 GND a_n55_n10# 0.21fF
C4 VDD w_15_7# 0.07fF
C5 GND B 0.16fF
C6 w_n28_13# out 0.06fF
C7 a_n55_n10# out 0.62fF
C8 a_n85_n22# w_n61_n20# 0.09fF
C9 B out 0.62fF
C10 a_n85_n22# VDD 0.41fF
C11 VDD A 0.19fF
C12 GND a_n85_n22# 0.21fF
C13 GND A 0.05fF
C14 a_n85_n22# out 0.12fF
C15 w_n98_8# a_n85_n22# 0.08fF
C16 w_n28_13# B 0.06fF
C17 a_n55_n10# B 0.07fF
C18 w_n98_8# A 0.09fF
C19 a_n55_n10# w_15_7# 0.08fF
C20 B w_15_7# 0.09fF
C21 out w_n61_n20# 0.06fF
C22 w_n28_13# A 0.09fF
C23 GND out 0.04fF
C24 a_n55_n10# A 0.40fF
C25 w_n98_8# VDD 0.07fF
C26 GND Gnd 1.25fF
C27 out Gnd 0.46fF
C28 a_n55_n10# Gnd 2.59fF
C29 B Gnd 0.03fF
C30 a_n85_n22# Gnd 1.72fF
C31 VDD Gnd 1.03fF
C32 A Gnd 3.13fF
C33 w_15_7# Gnd 1.43fF
C34 w_n28_13# Gnd 1.00fF
C35 w_n61_n20# Gnd 1.00fF
C36 w_n98_8# Gnd 1.43fF

    .tran 0.1n 200n
    .meas tran tpcq TRIG V(A) VAL=0.9 RISE=4
      + TARG V(out) VAL=0.9 FALL=1
    .control
    run
     set curplottitle  = "Eswar-2023102011"
    plot 6+v(A) 3+v(B) v(out)
    .endc
