magic
tech scmos
timestamp 1732375352
<< nwell >>
rect -735 75 -703 112
rect -697 75 -671 112
rect -653 75 -627 112
rect -608 75 -582 112
rect -522 75 -490 112
rect -484 75 -458 112
rect -440 75 -414 112
rect -395 75 -369 112
rect -275 25 -250 82
rect -238 -3 -213 37
rect -205 30 -180 70
rect -162 24 -137 81
rect -29 68 5 92
rect 11 67 35 91
rect 686 70 718 107
rect 724 70 750 107
rect 768 70 794 107
rect 813 70 839 107
rect 954 93 979 150
rect 991 65 1016 105
rect 1024 98 1049 138
rect 1067 92 1092 149
rect 1296 125 1328 162
rect 1334 125 1360 162
rect 1378 125 1404 162
rect 1423 125 1449 162
rect 254 -29 279 28
rect 291 -57 316 -17
rect 324 -24 349 16
rect 367 -30 392 27
rect 500 14 534 38
rect 540 13 564 37
rect 619 -34 653 2
rect 660 -35 684 -11
rect 505 -60 539 -36
rect 545 -61 569 -37
rect -720 -254 -688 -217
rect -682 -254 -656 -217
rect -638 -254 -612 -217
rect -593 -254 -567 -217
rect -507 -254 -475 -217
rect -469 -254 -443 -217
rect -425 -254 -399 -217
rect -380 -254 -354 -217
rect 249 -234 274 -177
rect -260 -304 -235 -247
rect -223 -332 -198 -292
rect -190 -299 -165 -259
rect -147 -305 -122 -248
rect -14 -261 20 -237
rect 26 -262 50 -238
rect 286 -262 311 -222
rect 319 -229 344 -189
rect 362 -235 387 -178
rect 495 -191 529 -167
rect 535 -192 559 -168
rect 614 -239 648 -203
rect 944 -215 969 -158
rect 655 -240 679 -216
rect 500 -265 534 -241
rect 540 -266 564 -242
rect 981 -243 1006 -203
rect 1014 -210 1039 -170
rect 1057 -216 1082 -159
rect 1286 -183 1318 -146
rect 1324 -183 1350 -146
rect 1368 -183 1394 -146
rect 1413 -183 1439 -146
rect -696 -521 -664 -484
rect -658 -521 -632 -484
rect -614 -521 -588 -484
rect -569 -521 -543 -484
rect -483 -521 -451 -484
rect -445 -521 -419 -484
rect -401 -521 -375 -484
rect -356 -521 -330 -484
rect 298 -488 323 -431
rect -236 -571 -211 -514
rect -199 -599 -174 -559
rect -166 -566 -141 -526
rect -123 -572 -98 -515
rect 10 -528 44 -504
rect 50 -529 74 -505
rect 335 -516 360 -476
rect 368 -483 393 -443
rect 411 -489 436 -432
rect 544 -445 578 -421
rect 584 -446 608 -422
rect 663 -493 697 -457
rect 704 -494 728 -470
rect 968 -474 993 -417
rect 549 -519 583 -495
rect 589 -520 613 -496
rect 1005 -502 1030 -462
rect 1038 -469 1063 -429
rect 1081 -475 1106 -418
rect 1310 -442 1342 -405
rect 1348 -442 1374 -405
rect 1392 -442 1418 -405
rect 1437 -442 1463 -405
rect 293 -693 318 -636
rect 330 -721 355 -681
rect 363 -688 388 -648
rect 406 -694 431 -637
rect 539 -650 573 -626
rect 579 -651 603 -627
rect 658 -698 692 -662
rect 699 -699 723 -675
rect 544 -724 578 -700
rect 584 -725 608 -701
rect 739 -708 771 -671
rect 777 -708 803 -671
rect 821 -708 847 -671
rect 866 -708 892 -671
rect 989 -780 1014 -723
rect -667 -831 -635 -794
rect -629 -831 -603 -794
rect -585 -831 -559 -794
rect -540 -831 -514 -794
rect -454 -831 -422 -794
rect -416 -831 -390 -794
rect -372 -831 -346 -794
rect -327 -831 -301 -794
rect 1026 -808 1051 -768
rect 1059 -775 1084 -735
rect 1102 -781 1127 -724
rect 1331 -748 1363 -711
rect 1369 -748 1395 -711
rect 1413 -748 1439 -711
rect 1458 -748 1484 -711
rect -207 -881 -182 -824
rect -170 -909 -145 -869
rect -137 -876 -112 -836
rect -94 -882 -69 -825
rect 39 -838 73 -814
rect 79 -839 103 -815
<< ntransistor >>
rect 1002 115 1004 135
rect -728 49 -726 59
rect -692 49 -690 59
rect -684 49 -682 59
rect -648 49 -646 59
rect -640 49 -638 59
rect -597 49 -595 59
rect -515 49 -513 59
rect -479 49 -477 59
rect -471 49 -469 59
rect -435 49 -433 59
rect -427 49 -425 59
rect -384 49 -382 59
rect -227 47 -225 67
rect -18 42 -16 54
rect -8 42 -6 54
rect 22 53 24 59
rect 965 63 967 83
rect 1035 68 1037 88
rect 1303 99 1305 109
rect 1339 99 1341 109
rect 1347 99 1349 109
rect 1383 99 1385 109
rect 1391 99 1393 109
rect 1434 99 1436 109
rect 1078 62 1080 82
rect 693 44 695 54
rect 729 44 731 54
rect 737 44 739 54
rect 773 44 775 54
rect 781 44 783 54
rect 824 44 826 54
rect -264 -5 -262 15
rect -194 0 -192 20
rect -151 -6 -149 14
rect 302 -7 304 13
rect 511 -12 513 0
rect 521 -12 523 0
rect 551 -1 553 5
rect 265 -59 267 -39
rect 335 -54 337 -34
rect 378 -60 380 -40
rect 671 -49 673 -43
rect 630 -55 632 -49
rect 640 -55 642 -49
rect 516 -86 518 -74
rect 526 -86 528 -74
rect 556 -75 558 -69
rect 297 -212 299 -192
rect -713 -280 -711 -270
rect -677 -280 -675 -270
rect -669 -280 -667 -270
rect -633 -280 -631 -270
rect -625 -280 -623 -270
rect -582 -280 -580 -270
rect -500 -280 -498 -270
rect -464 -280 -462 -270
rect -456 -280 -454 -270
rect -420 -280 -418 -270
rect -412 -280 -410 -270
rect -369 -280 -367 -270
rect 506 -217 508 -205
rect 516 -217 518 -205
rect 546 -206 548 -200
rect 992 -193 994 -173
rect -212 -282 -210 -262
rect 260 -264 262 -244
rect 330 -259 332 -239
rect 373 -265 375 -245
rect -3 -287 -1 -275
rect 7 -287 9 -275
rect 37 -276 39 -270
rect 955 -245 957 -225
rect 1025 -240 1027 -220
rect 1293 -209 1295 -199
rect 1329 -209 1331 -199
rect 1337 -209 1339 -199
rect 1373 -209 1375 -199
rect 1381 -209 1383 -199
rect 1424 -209 1426 -199
rect 1068 -246 1070 -226
rect 666 -254 668 -248
rect 625 -260 627 -254
rect 635 -260 637 -254
rect 511 -291 513 -279
rect 521 -291 523 -279
rect 551 -280 553 -274
rect -249 -334 -247 -314
rect -179 -329 -177 -309
rect -136 -335 -134 -315
rect 346 -466 348 -446
rect 555 -471 557 -459
rect 565 -471 567 -459
rect 595 -460 597 -454
rect -689 -547 -687 -537
rect -653 -547 -651 -537
rect -645 -547 -643 -537
rect -609 -547 -607 -537
rect -601 -547 -599 -537
rect -558 -547 -556 -537
rect -476 -547 -474 -537
rect -440 -547 -438 -537
rect -432 -547 -430 -537
rect -396 -547 -394 -537
rect -388 -547 -386 -537
rect -345 -547 -343 -537
rect -188 -549 -186 -529
rect 309 -518 311 -498
rect 379 -513 381 -493
rect 1016 -452 1018 -432
rect 422 -519 424 -499
rect 715 -508 717 -502
rect 979 -504 981 -484
rect 1049 -499 1051 -479
rect 1317 -468 1319 -458
rect 1353 -468 1355 -458
rect 1361 -468 1363 -458
rect 1397 -468 1399 -458
rect 1405 -468 1407 -458
rect 1448 -468 1450 -458
rect 1092 -505 1094 -485
rect 674 -514 676 -508
rect 684 -514 686 -508
rect 21 -554 23 -542
rect 31 -554 33 -542
rect 61 -543 63 -537
rect 560 -545 562 -533
rect 570 -545 572 -533
rect 600 -534 602 -528
rect -225 -601 -223 -581
rect -155 -596 -153 -576
rect -112 -602 -110 -582
rect 341 -671 343 -651
rect 550 -676 552 -664
rect 560 -676 562 -664
rect 590 -665 592 -659
rect 304 -723 306 -703
rect 374 -718 376 -698
rect 417 -724 419 -704
rect 710 -713 712 -707
rect 669 -719 671 -713
rect 679 -719 681 -713
rect 555 -750 557 -738
rect 565 -750 567 -738
rect 595 -739 597 -733
rect 746 -734 748 -724
rect 782 -734 784 -724
rect 790 -734 792 -724
rect 826 -734 828 -724
rect 834 -734 836 -724
rect 877 -734 879 -724
rect 1037 -758 1039 -738
rect 1000 -810 1002 -790
rect 1070 -805 1072 -785
rect 1338 -774 1340 -764
rect 1374 -774 1376 -764
rect 1382 -774 1384 -764
rect 1418 -774 1420 -764
rect 1426 -774 1428 -764
rect 1469 -774 1471 -764
rect 1113 -811 1115 -791
rect -660 -857 -658 -847
rect -624 -857 -622 -847
rect -616 -857 -614 -847
rect -580 -857 -578 -847
rect -572 -857 -570 -847
rect -529 -857 -527 -847
rect -447 -857 -445 -847
rect -411 -857 -409 -847
rect -403 -857 -401 -847
rect -367 -857 -365 -847
rect -359 -857 -357 -847
rect -316 -857 -314 -847
rect -159 -859 -157 -839
rect 50 -864 52 -852
rect 60 -864 62 -852
rect 90 -853 92 -847
rect -196 -911 -194 -891
rect -126 -906 -124 -886
rect -83 -912 -81 -892
<< ptransistor >>
rect -724 81 -722 106
rect -716 81 -714 106
rect -686 81 -684 106
rect -642 81 -640 106
rect -597 81 -595 106
rect -511 81 -509 106
rect -503 81 -501 106
rect -473 81 -471 106
rect -429 81 -427 106
rect -384 81 -382 106
rect 965 103 967 143
rect 1035 108 1037 128
rect -264 35 -262 75
rect -18 74 -16 86
rect -8 74 -6 86
rect -194 40 -192 60
rect -151 34 -149 74
rect 22 73 24 85
rect 697 76 699 101
rect 705 76 707 101
rect 735 76 737 101
rect 779 76 781 101
rect 824 76 826 101
rect 1078 102 1080 142
rect 1307 131 1309 156
rect 1315 131 1317 156
rect 1345 131 1347 156
rect 1389 131 1391 156
rect 1434 131 1436 156
rect 1002 75 1004 95
rect -227 7 -225 27
rect 265 -19 267 21
rect 511 20 513 32
rect 521 20 523 32
rect 335 -14 337 6
rect 378 -20 380 20
rect 551 19 553 31
rect 302 -47 304 -27
rect 630 -28 632 -4
rect 640 -28 642 -4
rect 516 -54 518 -42
rect 526 -54 528 -42
rect 556 -55 558 -43
rect 671 -29 673 -17
rect -709 -248 -707 -223
rect -701 -248 -699 -223
rect -671 -248 -669 -223
rect -627 -248 -625 -223
rect -582 -248 -580 -223
rect -496 -248 -494 -223
rect -488 -248 -486 -223
rect -458 -248 -456 -223
rect -414 -248 -412 -223
rect -369 -248 -367 -223
rect 260 -224 262 -184
rect 506 -185 508 -173
rect 516 -185 518 -173
rect 330 -219 332 -199
rect -249 -294 -247 -254
rect -3 -255 -1 -243
rect 7 -255 9 -243
rect 373 -225 375 -185
rect 546 -186 548 -174
rect 955 -205 957 -165
rect 1025 -200 1027 -180
rect -179 -289 -177 -269
rect -136 -295 -134 -255
rect 37 -256 39 -244
rect 297 -252 299 -232
rect 625 -233 627 -209
rect 635 -233 637 -209
rect 511 -259 513 -247
rect 521 -259 523 -247
rect 551 -260 553 -248
rect 666 -234 668 -222
rect 1068 -206 1070 -166
rect 1297 -177 1299 -152
rect 1305 -177 1307 -152
rect 1335 -177 1337 -152
rect 1379 -177 1381 -152
rect 1424 -177 1426 -152
rect 992 -233 994 -213
rect -212 -322 -210 -302
rect 309 -478 311 -438
rect 555 -439 557 -427
rect 565 -439 567 -427
rect 379 -473 381 -453
rect -685 -515 -683 -490
rect -677 -515 -675 -490
rect -647 -515 -645 -490
rect -603 -515 -601 -490
rect -558 -515 -556 -490
rect -472 -515 -470 -490
rect -464 -515 -462 -490
rect -434 -515 -432 -490
rect -390 -515 -388 -490
rect -345 -515 -343 -490
rect 422 -479 424 -439
rect 595 -440 597 -428
rect -225 -561 -223 -521
rect 21 -522 23 -510
rect 31 -522 33 -510
rect -155 -556 -153 -536
rect -112 -562 -110 -522
rect 61 -523 63 -511
rect 346 -506 348 -486
rect 674 -487 676 -463
rect 684 -487 686 -463
rect 979 -464 981 -424
rect 1049 -459 1051 -439
rect 560 -513 562 -501
rect 570 -513 572 -501
rect 600 -514 602 -502
rect 715 -488 717 -476
rect 1092 -465 1094 -425
rect 1321 -436 1323 -411
rect 1329 -436 1331 -411
rect 1359 -436 1361 -411
rect 1403 -436 1405 -411
rect 1448 -436 1450 -411
rect 1016 -492 1018 -472
rect -188 -589 -186 -569
rect 304 -683 306 -643
rect 550 -644 552 -632
rect 560 -644 562 -632
rect 374 -678 376 -658
rect 417 -684 419 -644
rect 590 -645 592 -633
rect 341 -711 343 -691
rect 669 -692 671 -668
rect 679 -692 681 -668
rect 555 -718 557 -706
rect 565 -718 567 -706
rect 595 -719 597 -707
rect 710 -693 712 -681
rect 750 -702 752 -677
rect 758 -702 760 -677
rect 788 -702 790 -677
rect 832 -702 834 -677
rect 877 -702 879 -677
rect 1000 -770 1002 -730
rect 1070 -765 1072 -745
rect 1113 -771 1115 -731
rect 1342 -742 1344 -717
rect 1350 -742 1352 -717
rect 1380 -742 1382 -717
rect 1424 -742 1426 -717
rect 1469 -742 1471 -717
rect -656 -825 -654 -800
rect -648 -825 -646 -800
rect -618 -825 -616 -800
rect -574 -825 -572 -800
rect -529 -825 -527 -800
rect -443 -825 -441 -800
rect -435 -825 -433 -800
rect -405 -825 -403 -800
rect -361 -825 -359 -800
rect -316 -825 -314 -800
rect 1037 -798 1039 -778
rect -196 -871 -194 -831
rect 50 -832 52 -820
rect 60 -832 62 -820
rect -126 -866 -124 -846
rect -83 -872 -81 -832
rect 90 -833 92 -821
rect -159 -899 -157 -879
<< ndiffusion >>
rect 1001 115 1002 135
rect 1004 115 1005 135
rect -729 49 -728 59
rect -726 49 -725 59
rect -693 49 -692 59
rect -690 49 -689 59
rect -685 49 -684 59
rect -682 49 -681 59
rect -649 49 -648 59
rect -646 49 -645 59
rect -641 49 -640 59
rect -638 49 -637 59
rect -598 49 -597 59
rect -595 49 -594 59
rect -516 49 -515 59
rect -513 49 -512 59
rect -480 49 -479 59
rect -477 49 -476 59
rect -472 49 -471 59
rect -469 49 -468 59
rect -436 49 -435 59
rect -433 49 -432 59
rect -428 49 -427 59
rect -425 49 -424 59
rect -385 49 -384 59
rect -382 49 -381 59
rect -228 47 -227 67
rect -225 47 -224 67
rect -19 42 -18 54
rect -16 42 -8 54
rect -6 42 -5 54
rect 21 53 22 59
rect 24 53 25 59
rect 964 63 965 83
rect 967 63 968 83
rect 1034 68 1035 88
rect 1037 68 1038 88
rect 1302 99 1303 109
rect 1305 99 1306 109
rect 1338 99 1339 109
rect 1341 99 1342 109
rect 1346 99 1347 109
rect 1349 99 1350 109
rect 1382 99 1383 109
rect 1385 99 1386 109
rect 1390 99 1391 109
rect 1393 99 1394 109
rect 1433 99 1434 109
rect 1436 99 1437 109
rect 1077 62 1078 82
rect 1080 62 1081 82
rect 692 44 693 54
rect 695 44 696 54
rect 728 44 729 54
rect 731 44 732 54
rect 736 44 737 54
rect 739 44 740 54
rect 772 44 773 54
rect 775 44 776 54
rect 780 44 781 54
rect 783 44 784 54
rect 823 44 824 54
rect 826 44 827 54
rect -265 -5 -264 15
rect -262 -5 -261 15
rect -195 0 -194 20
rect -192 0 -191 20
rect -152 -6 -151 14
rect -149 -6 -148 14
rect 301 -7 302 13
rect 304 -7 305 13
rect 510 -12 511 0
rect 513 -12 521 0
rect 523 -12 524 0
rect 550 -1 551 5
rect 553 -1 554 5
rect 264 -59 265 -39
rect 267 -59 268 -39
rect 334 -54 335 -34
rect 337 -54 338 -34
rect 377 -60 378 -40
rect 380 -60 381 -40
rect 670 -49 671 -43
rect 673 -49 674 -43
rect 629 -55 630 -49
rect 632 -55 634 -49
rect 638 -55 640 -49
rect 642 -55 643 -49
rect 515 -86 516 -74
rect 518 -86 526 -74
rect 528 -86 529 -74
rect 555 -75 556 -69
rect 558 -75 559 -69
rect 296 -212 297 -192
rect 299 -212 300 -192
rect -714 -280 -713 -270
rect -711 -280 -710 -270
rect -678 -280 -677 -270
rect -675 -280 -674 -270
rect -670 -280 -669 -270
rect -667 -280 -666 -270
rect -634 -280 -633 -270
rect -631 -280 -630 -270
rect -626 -280 -625 -270
rect -623 -280 -622 -270
rect -583 -280 -582 -270
rect -580 -280 -579 -270
rect -501 -280 -500 -270
rect -498 -280 -497 -270
rect -465 -280 -464 -270
rect -462 -280 -461 -270
rect -457 -280 -456 -270
rect -454 -280 -453 -270
rect -421 -280 -420 -270
rect -418 -280 -417 -270
rect -413 -280 -412 -270
rect -410 -280 -409 -270
rect -370 -280 -369 -270
rect -367 -280 -366 -270
rect 505 -217 506 -205
rect 508 -217 516 -205
rect 518 -217 519 -205
rect 545 -206 546 -200
rect 548 -206 549 -200
rect 991 -193 992 -173
rect 994 -193 995 -173
rect -213 -282 -212 -262
rect -210 -282 -209 -262
rect 259 -264 260 -244
rect 262 -264 263 -244
rect 329 -259 330 -239
rect 332 -259 333 -239
rect 372 -265 373 -245
rect 375 -265 376 -245
rect -4 -287 -3 -275
rect -1 -287 7 -275
rect 9 -287 10 -275
rect 36 -276 37 -270
rect 39 -276 40 -270
rect 954 -245 955 -225
rect 957 -245 958 -225
rect 1024 -240 1025 -220
rect 1027 -240 1028 -220
rect 1292 -209 1293 -199
rect 1295 -209 1296 -199
rect 1328 -209 1329 -199
rect 1331 -209 1332 -199
rect 1336 -209 1337 -199
rect 1339 -209 1340 -199
rect 1372 -209 1373 -199
rect 1375 -209 1376 -199
rect 1380 -209 1381 -199
rect 1383 -209 1384 -199
rect 1423 -209 1424 -199
rect 1426 -209 1427 -199
rect 1067 -246 1068 -226
rect 1070 -246 1071 -226
rect 665 -254 666 -248
rect 668 -254 669 -248
rect 624 -260 625 -254
rect 627 -260 629 -254
rect 633 -260 635 -254
rect 637 -260 638 -254
rect 510 -291 511 -279
rect 513 -291 521 -279
rect 523 -291 524 -279
rect 550 -280 551 -274
rect 553 -280 554 -274
rect -250 -334 -249 -314
rect -247 -334 -246 -314
rect -180 -329 -179 -309
rect -177 -329 -176 -309
rect -137 -335 -136 -315
rect -134 -335 -133 -315
rect 345 -466 346 -446
rect 348 -466 349 -446
rect 554 -471 555 -459
rect 557 -471 565 -459
rect 567 -471 568 -459
rect 594 -460 595 -454
rect 597 -460 598 -454
rect -690 -547 -689 -537
rect -687 -547 -686 -537
rect -654 -547 -653 -537
rect -651 -547 -650 -537
rect -646 -547 -645 -537
rect -643 -547 -642 -537
rect -610 -547 -609 -537
rect -607 -547 -606 -537
rect -602 -547 -601 -537
rect -599 -547 -598 -537
rect -559 -547 -558 -537
rect -556 -547 -555 -537
rect -477 -547 -476 -537
rect -474 -547 -473 -537
rect -441 -547 -440 -537
rect -438 -547 -437 -537
rect -433 -547 -432 -537
rect -430 -547 -429 -537
rect -397 -547 -396 -537
rect -394 -547 -393 -537
rect -389 -547 -388 -537
rect -386 -547 -385 -537
rect -346 -547 -345 -537
rect -343 -547 -342 -537
rect -189 -549 -188 -529
rect -186 -549 -185 -529
rect 308 -518 309 -498
rect 311 -518 312 -498
rect 378 -513 379 -493
rect 381 -513 382 -493
rect 1015 -452 1016 -432
rect 1018 -452 1019 -432
rect 421 -519 422 -499
rect 424 -519 425 -499
rect 714 -508 715 -502
rect 717 -508 718 -502
rect 978 -504 979 -484
rect 981 -504 982 -484
rect 1048 -499 1049 -479
rect 1051 -499 1052 -479
rect 1316 -468 1317 -458
rect 1319 -468 1320 -458
rect 1352 -468 1353 -458
rect 1355 -468 1356 -458
rect 1360 -468 1361 -458
rect 1363 -468 1364 -458
rect 1396 -468 1397 -458
rect 1399 -468 1400 -458
rect 1404 -468 1405 -458
rect 1407 -468 1408 -458
rect 1447 -468 1448 -458
rect 1450 -468 1451 -458
rect 1091 -505 1092 -485
rect 1094 -505 1095 -485
rect 673 -514 674 -508
rect 676 -514 678 -508
rect 682 -514 684 -508
rect 686 -514 687 -508
rect 20 -554 21 -542
rect 23 -554 31 -542
rect 33 -554 34 -542
rect 60 -543 61 -537
rect 63 -543 64 -537
rect 559 -545 560 -533
rect 562 -545 570 -533
rect 572 -545 573 -533
rect 599 -534 600 -528
rect 602 -534 603 -528
rect -226 -601 -225 -581
rect -223 -601 -222 -581
rect -156 -596 -155 -576
rect -153 -596 -152 -576
rect -113 -602 -112 -582
rect -110 -602 -109 -582
rect 340 -671 341 -651
rect 343 -671 344 -651
rect 549 -676 550 -664
rect 552 -676 560 -664
rect 562 -676 563 -664
rect 589 -665 590 -659
rect 592 -665 593 -659
rect 303 -723 304 -703
rect 306 -723 307 -703
rect 373 -718 374 -698
rect 376 -718 377 -698
rect 416 -724 417 -704
rect 419 -724 420 -704
rect 709 -713 710 -707
rect 712 -713 713 -707
rect 668 -719 669 -713
rect 671 -719 673 -713
rect 677 -719 679 -713
rect 681 -719 682 -713
rect 554 -750 555 -738
rect 557 -750 565 -738
rect 567 -750 568 -738
rect 594 -739 595 -733
rect 597 -739 598 -733
rect 745 -734 746 -724
rect 748 -734 749 -724
rect 781 -734 782 -724
rect 784 -734 785 -724
rect 789 -734 790 -724
rect 792 -734 793 -724
rect 825 -734 826 -724
rect 828 -734 829 -724
rect 833 -734 834 -724
rect 836 -734 837 -724
rect 876 -734 877 -724
rect 879 -734 880 -724
rect 1036 -758 1037 -738
rect 1039 -758 1040 -738
rect 999 -810 1000 -790
rect 1002 -810 1003 -790
rect 1069 -805 1070 -785
rect 1072 -805 1073 -785
rect 1337 -774 1338 -764
rect 1340 -774 1341 -764
rect 1373 -774 1374 -764
rect 1376 -774 1377 -764
rect 1381 -774 1382 -764
rect 1384 -774 1385 -764
rect 1417 -774 1418 -764
rect 1420 -774 1421 -764
rect 1425 -774 1426 -764
rect 1428 -774 1429 -764
rect 1468 -774 1469 -764
rect 1471 -774 1472 -764
rect 1112 -811 1113 -791
rect 1115 -811 1116 -791
rect -661 -857 -660 -847
rect -658 -857 -657 -847
rect -625 -857 -624 -847
rect -622 -857 -621 -847
rect -617 -857 -616 -847
rect -614 -857 -613 -847
rect -581 -857 -580 -847
rect -578 -857 -577 -847
rect -573 -857 -572 -847
rect -570 -857 -569 -847
rect -530 -857 -529 -847
rect -527 -857 -526 -847
rect -448 -857 -447 -847
rect -445 -857 -444 -847
rect -412 -857 -411 -847
rect -409 -857 -408 -847
rect -404 -857 -403 -847
rect -401 -857 -400 -847
rect -368 -857 -367 -847
rect -365 -857 -364 -847
rect -360 -857 -359 -847
rect -357 -857 -356 -847
rect -317 -857 -316 -847
rect -314 -857 -313 -847
rect -160 -859 -159 -839
rect -157 -859 -156 -839
rect 49 -864 50 -852
rect 52 -864 60 -852
rect 62 -864 63 -852
rect 89 -853 90 -847
rect 92 -853 93 -847
rect -197 -911 -196 -891
rect -194 -911 -193 -891
rect -127 -906 -126 -886
rect -124 -906 -123 -886
rect -84 -912 -83 -892
rect -81 -912 -80 -892
<< pdiffusion >>
rect -725 81 -724 106
rect -722 81 -721 106
rect -717 81 -716 106
rect -714 81 -713 106
rect -687 81 -686 106
rect -684 81 -683 106
rect -643 81 -642 106
rect -640 81 -639 106
rect -598 81 -597 106
rect -595 81 -594 106
rect -512 81 -511 106
rect -509 81 -508 106
rect -504 81 -503 106
rect -501 81 -500 106
rect -474 81 -473 106
rect -471 81 -470 106
rect -430 81 -429 106
rect -427 81 -426 106
rect -385 81 -384 106
rect -382 81 -381 106
rect 964 103 965 143
rect 967 103 968 143
rect 1034 108 1035 128
rect 1037 108 1038 128
rect -265 35 -264 75
rect -262 35 -261 75
rect -19 74 -18 86
rect -16 74 -14 86
rect -10 74 -8 86
rect -6 74 -5 86
rect -195 40 -194 60
rect -192 40 -191 60
rect -152 34 -151 74
rect -149 34 -148 74
rect 21 73 22 85
rect 24 73 25 85
rect 696 76 697 101
rect 699 76 700 101
rect 704 76 705 101
rect 707 76 708 101
rect 734 76 735 101
rect 737 76 738 101
rect 778 76 779 101
rect 781 76 782 101
rect 823 76 824 101
rect 826 76 827 101
rect 1077 102 1078 142
rect 1080 102 1081 142
rect 1306 131 1307 156
rect 1309 131 1310 156
rect 1314 131 1315 156
rect 1317 131 1318 156
rect 1344 131 1345 156
rect 1347 131 1348 156
rect 1388 131 1389 156
rect 1391 131 1392 156
rect 1433 131 1434 156
rect 1436 131 1437 156
rect 1001 75 1002 95
rect 1004 75 1005 95
rect -228 7 -227 27
rect -225 7 -224 27
rect 264 -19 265 21
rect 267 -19 268 21
rect 510 20 511 32
rect 513 20 515 32
rect 519 20 521 32
rect 523 20 524 32
rect 334 -14 335 6
rect 337 -14 338 6
rect 377 -20 378 20
rect 380 -20 381 20
rect 550 19 551 31
rect 553 19 554 31
rect 301 -47 302 -27
rect 304 -47 305 -27
rect 629 -28 630 -4
rect 632 -28 640 -4
rect 642 -28 643 -4
rect 515 -54 516 -42
rect 518 -54 520 -42
rect 524 -54 526 -42
rect 528 -54 529 -42
rect 555 -55 556 -43
rect 558 -55 559 -43
rect 670 -29 671 -17
rect 673 -29 674 -17
rect -710 -248 -709 -223
rect -707 -248 -706 -223
rect -702 -248 -701 -223
rect -699 -248 -698 -223
rect -672 -248 -671 -223
rect -669 -248 -668 -223
rect -628 -248 -627 -223
rect -625 -248 -624 -223
rect -583 -248 -582 -223
rect -580 -248 -579 -223
rect -497 -248 -496 -223
rect -494 -248 -493 -223
rect -489 -248 -488 -223
rect -486 -248 -485 -223
rect -459 -248 -458 -223
rect -456 -248 -455 -223
rect -415 -248 -414 -223
rect -412 -248 -411 -223
rect -370 -248 -369 -223
rect -367 -248 -366 -223
rect 259 -224 260 -184
rect 262 -224 263 -184
rect 505 -185 506 -173
rect 508 -185 510 -173
rect 514 -185 516 -173
rect 518 -185 519 -173
rect 329 -219 330 -199
rect 332 -219 333 -199
rect -250 -294 -249 -254
rect -247 -294 -246 -254
rect -4 -255 -3 -243
rect -1 -255 1 -243
rect 5 -255 7 -243
rect 9 -255 10 -243
rect 372 -225 373 -185
rect 375 -225 376 -185
rect 545 -186 546 -174
rect 548 -186 549 -174
rect 954 -205 955 -165
rect 957 -205 958 -165
rect 1024 -200 1025 -180
rect 1027 -200 1028 -180
rect -180 -289 -179 -269
rect -177 -289 -176 -269
rect -137 -295 -136 -255
rect -134 -295 -133 -255
rect 36 -256 37 -244
rect 39 -256 40 -244
rect 296 -252 297 -232
rect 299 -252 300 -232
rect 624 -233 625 -209
rect 627 -233 635 -209
rect 637 -233 638 -209
rect 510 -259 511 -247
rect 513 -259 515 -247
rect 519 -259 521 -247
rect 523 -259 524 -247
rect 550 -260 551 -248
rect 553 -260 554 -248
rect 665 -234 666 -222
rect 668 -234 669 -222
rect 1067 -206 1068 -166
rect 1070 -206 1071 -166
rect 1296 -177 1297 -152
rect 1299 -177 1300 -152
rect 1304 -177 1305 -152
rect 1307 -177 1308 -152
rect 1334 -177 1335 -152
rect 1337 -177 1338 -152
rect 1378 -177 1379 -152
rect 1381 -177 1382 -152
rect 1423 -177 1424 -152
rect 1426 -177 1427 -152
rect 991 -233 992 -213
rect 994 -233 995 -213
rect -213 -322 -212 -302
rect -210 -322 -209 -302
rect 308 -478 309 -438
rect 311 -478 312 -438
rect 554 -439 555 -427
rect 557 -439 559 -427
rect 563 -439 565 -427
rect 567 -439 568 -427
rect 378 -473 379 -453
rect 381 -473 382 -453
rect -686 -515 -685 -490
rect -683 -515 -682 -490
rect -678 -515 -677 -490
rect -675 -515 -674 -490
rect -648 -515 -647 -490
rect -645 -515 -644 -490
rect -604 -515 -603 -490
rect -601 -515 -600 -490
rect -559 -515 -558 -490
rect -556 -515 -555 -490
rect -473 -515 -472 -490
rect -470 -515 -469 -490
rect -465 -515 -464 -490
rect -462 -515 -461 -490
rect -435 -515 -434 -490
rect -432 -515 -431 -490
rect -391 -515 -390 -490
rect -388 -515 -387 -490
rect -346 -515 -345 -490
rect -343 -515 -342 -490
rect 421 -479 422 -439
rect 424 -479 425 -439
rect 594 -440 595 -428
rect 597 -440 598 -428
rect -226 -561 -225 -521
rect -223 -561 -222 -521
rect 20 -522 21 -510
rect 23 -522 25 -510
rect 29 -522 31 -510
rect 33 -522 34 -510
rect -156 -556 -155 -536
rect -153 -556 -152 -536
rect -113 -562 -112 -522
rect -110 -562 -109 -522
rect 60 -523 61 -511
rect 63 -523 64 -511
rect 345 -506 346 -486
rect 348 -506 349 -486
rect 673 -487 674 -463
rect 676 -487 684 -463
rect 686 -487 687 -463
rect 978 -464 979 -424
rect 981 -464 982 -424
rect 1048 -459 1049 -439
rect 1051 -459 1052 -439
rect 559 -513 560 -501
rect 562 -513 564 -501
rect 568 -513 570 -501
rect 572 -513 573 -501
rect 599 -514 600 -502
rect 602 -514 603 -502
rect 714 -488 715 -476
rect 717 -488 718 -476
rect 1091 -465 1092 -425
rect 1094 -465 1095 -425
rect 1320 -436 1321 -411
rect 1323 -436 1324 -411
rect 1328 -436 1329 -411
rect 1331 -436 1332 -411
rect 1358 -436 1359 -411
rect 1361 -436 1362 -411
rect 1402 -436 1403 -411
rect 1405 -436 1406 -411
rect 1447 -436 1448 -411
rect 1450 -436 1451 -411
rect 1015 -492 1016 -472
rect 1018 -492 1019 -472
rect -189 -589 -188 -569
rect -186 -589 -185 -569
rect 303 -683 304 -643
rect 306 -683 307 -643
rect 549 -644 550 -632
rect 552 -644 554 -632
rect 558 -644 560 -632
rect 562 -644 563 -632
rect 373 -678 374 -658
rect 376 -678 377 -658
rect 416 -684 417 -644
rect 419 -684 420 -644
rect 589 -645 590 -633
rect 592 -645 593 -633
rect 340 -711 341 -691
rect 343 -711 344 -691
rect 668 -692 669 -668
rect 671 -692 679 -668
rect 681 -692 682 -668
rect 554 -718 555 -706
rect 557 -718 559 -706
rect 563 -718 565 -706
rect 567 -718 568 -706
rect 594 -719 595 -707
rect 597 -719 598 -707
rect 709 -693 710 -681
rect 712 -693 713 -681
rect 749 -702 750 -677
rect 752 -702 753 -677
rect 757 -702 758 -677
rect 760 -702 761 -677
rect 787 -702 788 -677
rect 790 -702 791 -677
rect 831 -702 832 -677
rect 834 -702 835 -677
rect 876 -702 877 -677
rect 879 -702 880 -677
rect 999 -770 1000 -730
rect 1002 -770 1003 -730
rect 1069 -765 1070 -745
rect 1072 -765 1073 -745
rect 1112 -771 1113 -731
rect 1115 -771 1116 -731
rect 1341 -742 1342 -717
rect 1344 -742 1345 -717
rect 1349 -742 1350 -717
rect 1352 -742 1353 -717
rect 1379 -742 1380 -717
rect 1382 -742 1383 -717
rect 1423 -742 1424 -717
rect 1426 -742 1427 -717
rect 1468 -742 1469 -717
rect 1471 -742 1472 -717
rect -657 -825 -656 -800
rect -654 -825 -653 -800
rect -649 -825 -648 -800
rect -646 -825 -645 -800
rect -619 -825 -618 -800
rect -616 -825 -615 -800
rect -575 -825 -574 -800
rect -572 -825 -571 -800
rect -530 -825 -529 -800
rect -527 -825 -526 -800
rect -444 -825 -443 -800
rect -441 -825 -440 -800
rect -436 -825 -435 -800
rect -433 -825 -432 -800
rect -406 -825 -405 -800
rect -403 -825 -402 -800
rect -362 -825 -361 -800
rect -359 -825 -358 -800
rect -317 -825 -316 -800
rect -314 -825 -313 -800
rect 1036 -798 1037 -778
rect 1039 -798 1040 -778
rect -197 -871 -196 -831
rect -194 -871 -193 -831
rect 49 -832 50 -820
rect 52 -832 54 -820
rect 58 -832 60 -820
rect 62 -832 63 -820
rect -127 -866 -126 -846
rect -124 -866 -123 -846
rect -84 -872 -83 -832
rect -81 -872 -80 -832
rect 89 -833 90 -821
rect 92 -833 93 -821
rect -160 -899 -159 -879
rect -157 -899 -156 -879
<< ndcontact >>
rect 997 115 1001 135
rect 1005 115 1009 135
rect -733 49 -729 59
rect -725 49 -721 59
rect -697 49 -693 59
rect -689 49 -685 59
rect -681 49 -677 59
rect -653 49 -649 59
rect -645 49 -641 59
rect -637 49 -633 59
rect -602 49 -598 59
rect -594 49 -590 59
rect -520 49 -516 59
rect -512 49 -508 59
rect -484 49 -480 59
rect -476 49 -472 59
rect -468 49 -464 59
rect -440 49 -436 59
rect -432 49 -428 59
rect -424 49 -420 59
rect -389 49 -385 59
rect -381 49 -377 59
rect -232 47 -228 67
rect -224 47 -220 67
rect -23 42 -19 54
rect -5 42 -1 54
rect 17 53 21 59
rect 25 53 29 59
rect 960 63 964 83
rect 968 63 972 83
rect 1030 68 1034 88
rect 1038 68 1042 88
rect 1298 99 1302 109
rect 1306 99 1310 109
rect 1334 99 1338 109
rect 1342 99 1346 109
rect 1350 99 1354 109
rect 1378 99 1382 109
rect 1386 99 1390 109
rect 1394 99 1398 109
rect 1429 99 1433 109
rect 1437 99 1441 109
rect 1073 62 1077 82
rect 1081 62 1085 82
rect 688 44 692 54
rect 696 44 700 54
rect 724 44 728 54
rect 732 44 736 54
rect 740 44 744 54
rect 768 44 772 54
rect 776 44 780 54
rect 784 44 788 54
rect 819 44 823 54
rect 827 44 831 54
rect -269 -5 -265 15
rect -261 -5 -257 15
rect -199 0 -195 20
rect -191 0 -187 20
rect -156 -6 -152 14
rect -148 -6 -144 14
rect 297 -7 301 13
rect 305 -7 309 13
rect 506 -12 510 0
rect 524 -12 528 0
rect 546 -1 550 5
rect 554 -1 558 5
rect 260 -59 264 -39
rect 268 -59 272 -39
rect 330 -54 334 -34
rect 338 -54 342 -34
rect 373 -60 377 -40
rect 381 -60 385 -40
rect 666 -49 670 -43
rect 674 -49 678 -43
rect 625 -55 629 -49
rect 634 -55 638 -49
rect 643 -55 647 -49
rect 511 -86 515 -74
rect 529 -86 533 -74
rect 551 -75 555 -69
rect 559 -75 563 -69
rect 292 -212 296 -192
rect 300 -212 304 -192
rect -718 -280 -714 -270
rect -710 -280 -706 -270
rect -682 -280 -678 -270
rect -674 -280 -670 -270
rect -666 -280 -662 -270
rect -638 -280 -634 -270
rect -630 -280 -626 -270
rect -622 -280 -618 -270
rect -587 -280 -583 -270
rect -579 -280 -575 -270
rect -505 -280 -501 -270
rect -497 -280 -493 -270
rect -469 -280 -465 -270
rect -461 -280 -457 -270
rect -453 -280 -449 -270
rect -425 -280 -421 -270
rect -417 -280 -413 -270
rect -409 -280 -405 -270
rect -374 -280 -370 -270
rect -366 -280 -362 -270
rect 501 -217 505 -205
rect 519 -217 523 -205
rect 541 -206 545 -200
rect 549 -206 553 -200
rect 987 -193 991 -173
rect 995 -193 999 -173
rect -217 -282 -213 -262
rect -209 -282 -205 -262
rect 255 -264 259 -244
rect 263 -264 267 -244
rect 325 -259 329 -239
rect 333 -259 337 -239
rect 368 -265 372 -245
rect 376 -265 380 -245
rect -8 -287 -4 -275
rect 10 -287 14 -275
rect 32 -276 36 -270
rect 40 -276 44 -270
rect 950 -245 954 -225
rect 958 -245 962 -225
rect 1020 -240 1024 -220
rect 1028 -240 1032 -220
rect 1288 -209 1292 -199
rect 1296 -209 1300 -199
rect 1324 -209 1328 -199
rect 1332 -209 1336 -199
rect 1340 -209 1344 -199
rect 1368 -209 1372 -199
rect 1376 -209 1380 -199
rect 1384 -209 1388 -199
rect 1419 -209 1423 -199
rect 1427 -209 1431 -199
rect 1063 -246 1067 -226
rect 1071 -246 1075 -226
rect 661 -254 665 -248
rect 669 -254 673 -248
rect 620 -260 624 -254
rect 629 -260 633 -254
rect 638 -260 642 -254
rect 506 -291 510 -279
rect 524 -291 528 -279
rect 546 -280 550 -274
rect 554 -280 558 -274
rect -254 -334 -250 -314
rect -246 -334 -242 -314
rect -184 -329 -180 -309
rect -176 -329 -172 -309
rect -141 -335 -137 -315
rect -133 -335 -129 -315
rect 341 -466 345 -446
rect 349 -466 353 -446
rect 550 -471 554 -459
rect 568 -471 572 -459
rect 590 -460 594 -454
rect 598 -460 602 -454
rect -694 -547 -690 -537
rect -686 -547 -682 -537
rect -658 -547 -654 -537
rect -650 -547 -646 -537
rect -642 -547 -638 -537
rect -614 -547 -610 -537
rect -606 -547 -602 -537
rect -598 -547 -594 -537
rect -563 -547 -559 -537
rect -555 -547 -551 -537
rect -481 -547 -477 -537
rect -473 -547 -469 -537
rect -445 -547 -441 -537
rect -437 -547 -433 -537
rect -429 -547 -425 -537
rect -401 -547 -397 -537
rect -393 -547 -389 -537
rect -385 -547 -381 -537
rect -350 -547 -346 -537
rect -342 -547 -338 -537
rect -193 -549 -189 -529
rect -185 -549 -181 -529
rect 304 -518 308 -498
rect 312 -518 316 -498
rect 374 -513 378 -493
rect 382 -513 386 -493
rect 1011 -452 1015 -432
rect 1019 -452 1023 -432
rect 417 -519 421 -499
rect 425 -519 429 -499
rect 710 -508 714 -502
rect 718 -508 722 -502
rect 974 -504 978 -484
rect 982 -504 986 -484
rect 1044 -499 1048 -479
rect 1052 -499 1056 -479
rect 1312 -468 1316 -458
rect 1320 -468 1324 -458
rect 1348 -468 1352 -458
rect 1356 -468 1360 -458
rect 1364 -468 1368 -458
rect 1392 -468 1396 -458
rect 1400 -468 1404 -458
rect 1408 -468 1412 -458
rect 1443 -468 1447 -458
rect 1451 -468 1455 -458
rect 1087 -505 1091 -485
rect 1095 -505 1099 -485
rect 669 -514 673 -508
rect 678 -514 682 -508
rect 687 -514 691 -508
rect 16 -554 20 -542
rect 34 -554 38 -542
rect 56 -543 60 -537
rect 64 -543 68 -537
rect 555 -545 559 -533
rect 573 -545 577 -533
rect 595 -534 599 -528
rect 603 -534 607 -528
rect -230 -601 -226 -581
rect -222 -601 -218 -581
rect -160 -596 -156 -576
rect -152 -596 -148 -576
rect -117 -602 -113 -582
rect -109 -602 -105 -582
rect 336 -671 340 -651
rect 344 -671 348 -651
rect 545 -676 549 -664
rect 563 -676 567 -664
rect 585 -665 589 -659
rect 593 -665 597 -659
rect 299 -723 303 -703
rect 307 -723 311 -703
rect 369 -718 373 -698
rect 377 -718 381 -698
rect 412 -724 416 -704
rect 420 -724 424 -704
rect 705 -713 709 -707
rect 713 -713 717 -707
rect 664 -719 668 -713
rect 673 -719 677 -713
rect 682 -719 686 -713
rect 550 -750 554 -738
rect 568 -750 572 -738
rect 590 -739 594 -733
rect 598 -739 602 -733
rect 741 -734 745 -724
rect 749 -734 753 -724
rect 777 -734 781 -724
rect 785 -734 789 -724
rect 793 -734 797 -724
rect 821 -734 825 -724
rect 829 -734 833 -724
rect 837 -734 841 -724
rect 872 -734 876 -724
rect 880 -734 884 -724
rect 1032 -758 1036 -738
rect 1040 -758 1044 -738
rect 995 -810 999 -790
rect 1003 -810 1007 -790
rect 1065 -805 1069 -785
rect 1073 -805 1077 -785
rect 1333 -774 1337 -764
rect 1341 -774 1345 -764
rect 1369 -774 1373 -764
rect 1377 -774 1381 -764
rect 1385 -774 1389 -764
rect 1413 -774 1417 -764
rect 1421 -774 1425 -764
rect 1429 -774 1433 -764
rect 1464 -774 1468 -764
rect 1472 -774 1476 -764
rect 1108 -811 1112 -791
rect 1116 -811 1120 -791
rect -665 -857 -661 -847
rect -657 -857 -653 -847
rect -629 -857 -625 -847
rect -621 -857 -617 -847
rect -613 -857 -609 -847
rect -585 -857 -581 -847
rect -577 -857 -573 -847
rect -569 -857 -565 -847
rect -534 -857 -530 -847
rect -526 -857 -522 -847
rect -452 -857 -448 -847
rect -444 -857 -440 -847
rect -416 -857 -412 -847
rect -408 -857 -404 -847
rect -400 -857 -396 -847
rect -372 -857 -368 -847
rect -364 -857 -360 -847
rect -356 -857 -352 -847
rect -321 -857 -317 -847
rect -313 -857 -309 -847
rect -164 -859 -160 -839
rect -156 -859 -152 -839
rect 45 -864 49 -852
rect 63 -864 67 -852
rect 85 -853 89 -847
rect 93 -853 97 -847
rect -201 -911 -197 -891
rect -193 -911 -189 -891
rect -131 -906 -127 -886
rect -123 -906 -119 -886
rect -88 -912 -84 -892
rect -80 -912 -76 -892
<< pdcontact >>
rect -729 81 -725 106
rect -721 81 -717 106
rect -713 81 -709 106
rect -691 81 -687 106
rect -683 81 -679 106
rect -647 81 -643 106
rect -639 81 -635 106
rect -602 81 -598 106
rect -594 81 -590 106
rect -516 81 -512 106
rect -508 81 -504 106
rect -500 81 -496 106
rect -478 81 -474 106
rect -470 81 -466 106
rect -434 81 -430 106
rect -426 81 -422 106
rect -389 81 -385 106
rect -381 81 -377 106
rect 960 103 964 143
rect 968 103 972 143
rect 1030 108 1034 128
rect 1038 108 1042 128
rect -269 35 -265 75
rect -261 35 -257 75
rect -23 74 -19 86
rect -14 74 -10 86
rect -5 74 -1 86
rect -199 40 -195 60
rect -191 40 -187 60
rect -156 34 -152 74
rect -148 34 -144 74
rect 17 73 21 85
rect 25 73 29 85
rect 692 76 696 101
rect 700 76 704 101
rect 708 76 712 101
rect 730 76 734 101
rect 738 76 742 101
rect 774 76 778 101
rect 782 76 786 101
rect 819 76 823 101
rect 827 76 831 101
rect 1073 102 1077 142
rect 1081 102 1085 142
rect 1302 131 1306 156
rect 1310 131 1314 156
rect 1318 131 1322 156
rect 1340 131 1344 156
rect 1348 131 1352 156
rect 1384 131 1388 156
rect 1392 131 1396 156
rect 1429 131 1433 156
rect 1437 131 1441 156
rect 997 75 1001 95
rect 1005 75 1009 95
rect -232 7 -228 27
rect -224 7 -220 27
rect 260 -19 264 21
rect 268 -19 272 21
rect 506 20 510 32
rect 515 20 519 32
rect 524 20 528 32
rect 330 -14 334 6
rect 338 -14 342 6
rect 373 -20 377 20
rect 381 -20 385 20
rect 546 19 550 31
rect 554 19 558 31
rect 297 -47 301 -27
rect 305 -47 309 -27
rect 625 -28 629 -4
rect 643 -28 647 -4
rect 511 -54 515 -42
rect 520 -54 524 -42
rect 529 -54 533 -42
rect 551 -55 555 -43
rect 559 -55 563 -43
rect 666 -29 670 -17
rect 674 -29 678 -17
rect -714 -248 -710 -223
rect -706 -248 -702 -223
rect -698 -248 -694 -223
rect -676 -248 -672 -223
rect -668 -248 -664 -223
rect -632 -248 -628 -223
rect -624 -248 -620 -223
rect -587 -248 -583 -223
rect -579 -248 -575 -223
rect -501 -248 -497 -223
rect -493 -248 -489 -223
rect -485 -248 -481 -223
rect -463 -248 -459 -223
rect -455 -248 -451 -223
rect -419 -248 -415 -223
rect -411 -248 -407 -223
rect -374 -248 -370 -223
rect -366 -248 -362 -223
rect 255 -224 259 -184
rect 263 -224 267 -184
rect 501 -185 505 -173
rect 510 -185 514 -173
rect 519 -185 523 -173
rect 325 -219 329 -199
rect 333 -219 337 -199
rect -254 -294 -250 -254
rect -246 -294 -242 -254
rect -8 -255 -4 -243
rect 1 -255 5 -243
rect 10 -255 14 -243
rect 368 -225 372 -185
rect 376 -225 380 -185
rect 541 -186 545 -174
rect 549 -186 553 -174
rect 950 -205 954 -165
rect 958 -205 962 -165
rect 1020 -200 1024 -180
rect 1028 -200 1032 -180
rect -184 -289 -180 -269
rect -176 -289 -172 -269
rect -141 -295 -137 -255
rect -133 -295 -129 -255
rect 32 -256 36 -244
rect 40 -256 44 -244
rect 292 -252 296 -232
rect 300 -252 304 -232
rect 620 -233 624 -209
rect 638 -233 642 -209
rect 506 -259 510 -247
rect 515 -259 519 -247
rect 524 -259 528 -247
rect 546 -260 550 -248
rect 554 -260 558 -248
rect 661 -234 665 -222
rect 669 -234 673 -222
rect 1063 -206 1067 -166
rect 1071 -206 1075 -166
rect 1292 -177 1296 -152
rect 1300 -177 1304 -152
rect 1308 -177 1312 -152
rect 1330 -177 1334 -152
rect 1338 -177 1342 -152
rect 1374 -177 1378 -152
rect 1382 -177 1386 -152
rect 1419 -177 1423 -152
rect 1427 -177 1431 -152
rect 987 -233 991 -213
rect 995 -233 999 -213
rect -217 -322 -213 -302
rect -209 -322 -205 -302
rect 304 -478 308 -438
rect 312 -478 316 -438
rect 550 -439 554 -427
rect 559 -439 563 -427
rect 568 -439 572 -427
rect 374 -473 378 -453
rect 382 -473 386 -453
rect -690 -515 -686 -490
rect -682 -515 -678 -490
rect -674 -515 -670 -490
rect -652 -515 -648 -490
rect -644 -515 -640 -490
rect -608 -515 -604 -490
rect -600 -515 -596 -490
rect -563 -515 -559 -490
rect -555 -515 -551 -490
rect -477 -515 -473 -490
rect -469 -515 -465 -490
rect -461 -515 -457 -490
rect -439 -515 -435 -490
rect -431 -515 -427 -490
rect -395 -515 -391 -490
rect -387 -515 -383 -490
rect -350 -515 -346 -490
rect -342 -515 -338 -490
rect 417 -479 421 -439
rect 425 -479 429 -439
rect 590 -440 594 -428
rect 598 -440 602 -428
rect -230 -561 -226 -521
rect -222 -561 -218 -521
rect 16 -522 20 -510
rect 25 -522 29 -510
rect 34 -522 38 -510
rect -160 -556 -156 -536
rect -152 -556 -148 -536
rect -117 -562 -113 -522
rect -109 -562 -105 -522
rect 56 -523 60 -511
rect 64 -523 68 -511
rect 341 -506 345 -486
rect 349 -506 353 -486
rect 669 -487 673 -463
rect 687 -487 691 -463
rect 974 -464 978 -424
rect 982 -464 986 -424
rect 1044 -459 1048 -439
rect 1052 -459 1056 -439
rect 555 -513 559 -501
rect 564 -513 568 -501
rect 573 -513 577 -501
rect 595 -514 599 -502
rect 603 -514 607 -502
rect 710 -488 714 -476
rect 718 -488 722 -476
rect 1087 -465 1091 -425
rect 1095 -465 1099 -425
rect 1316 -436 1320 -411
rect 1324 -436 1328 -411
rect 1332 -436 1336 -411
rect 1354 -436 1358 -411
rect 1362 -436 1366 -411
rect 1398 -436 1402 -411
rect 1406 -436 1410 -411
rect 1443 -436 1447 -411
rect 1451 -436 1455 -411
rect 1011 -492 1015 -472
rect 1019 -492 1023 -472
rect -193 -589 -189 -569
rect -185 -589 -181 -569
rect 299 -683 303 -643
rect 307 -683 311 -643
rect 545 -644 549 -632
rect 554 -644 558 -632
rect 563 -644 567 -632
rect 369 -678 373 -658
rect 377 -678 381 -658
rect 412 -684 416 -644
rect 420 -684 424 -644
rect 585 -645 589 -633
rect 593 -645 597 -633
rect 336 -711 340 -691
rect 344 -711 348 -691
rect 664 -692 668 -668
rect 682 -692 686 -668
rect 550 -718 554 -706
rect 559 -718 563 -706
rect 568 -718 572 -706
rect 590 -719 594 -707
rect 598 -719 602 -707
rect 705 -693 709 -681
rect 713 -693 717 -681
rect 745 -702 749 -677
rect 753 -702 757 -677
rect 761 -702 765 -677
rect 783 -702 787 -677
rect 791 -702 795 -677
rect 827 -702 831 -677
rect 835 -702 839 -677
rect 872 -702 876 -677
rect 880 -702 884 -677
rect 995 -770 999 -730
rect 1003 -770 1007 -730
rect 1065 -765 1069 -745
rect 1073 -765 1077 -745
rect 1108 -771 1112 -731
rect 1116 -771 1120 -731
rect 1337 -742 1341 -717
rect 1345 -742 1349 -717
rect 1353 -742 1357 -717
rect 1375 -742 1379 -717
rect 1383 -742 1387 -717
rect 1419 -742 1423 -717
rect 1427 -742 1431 -717
rect 1464 -742 1468 -717
rect 1472 -742 1476 -717
rect -661 -825 -657 -800
rect -653 -825 -649 -800
rect -645 -825 -641 -800
rect -623 -825 -619 -800
rect -615 -825 -611 -800
rect -579 -825 -575 -800
rect -571 -825 -567 -800
rect -534 -825 -530 -800
rect -526 -825 -522 -800
rect -448 -825 -444 -800
rect -440 -825 -436 -800
rect -432 -825 -428 -800
rect -410 -825 -406 -800
rect -402 -825 -398 -800
rect -366 -825 -362 -800
rect -358 -825 -354 -800
rect -321 -825 -317 -800
rect -313 -825 -309 -800
rect 1032 -798 1036 -778
rect 1040 -798 1044 -778
rect -201 -871 -197 -831
rect -193 -871 -189 -831
rect 45 -832 49 -820
rect 54 -832 58 -820
rect 63 -832 67 -820
rect -131 -866 -127 -846
rect -123 -866 -119 -846
rect -88 -872 -84 -832
rect -80 -872 -76 -832
rect 85 -833 89 -821
rect 93 -833 97 -821
rect -164 -899 -160 -879
rect -156 -899 -152 -879
<< polysilicon >>
rect 1307 156 1309 159
rect 1315 156 1317 159
rect 1345 156 1347 159
rect 1389 156 1391 159
rect 1434 156 1436 159
rect 965 143 967 147
rect -724 106 -722 109
rect -716 106 -714 109
rect -686 106 -684 109
rect -642 106 -640 109
rect -597 106 -595 109
rect -511 106 -509 109
rect -503 106 -501 109
rect -473 106 -471 109
rect -429 106 -427 109
rect -384 106 -382 109
rect 697 101 699 104
rect 705 101 707 104
rect 735 101 737 104
rect 779 101 781 104
rect 824 101 826 104
rect 1078 142 1080 146
rect 1002 135 1004 142
rect 1035 128 1037 142
rect 1002 112 1004 115
rect 1035 105 1037 108
rect -18 86 -16 89
rect -8 86 -6 89
rect -724 74 -722 81
rect -729 70 -722 74
rect -728 59 -726 70
rect -716 62 -714 81
rect -686 73 -684 81
rect -642 73 -640 81
rect -692 71 -684 73
rect -648 71 -640 73
rect -692 59 -690 71
rect -684 59 -682 68
rect -648 59 -646 71
rect -640 59 -638 68
rect -597 59 -595 81
rect -511 74 -509 81
rect -516 70 -509 74
rect -515 59 -513 70
rect -503 62 -501 81
rect -473 73 -471 81
rect -429 73 -427 81
rect -479 71 -471 73
rect -435 71 -427 73
rect -479 59 -477 71
rect -471 59 -469 68
rect -435 59 -433 71
rect -427 59 -425 68
rect -384 59 -382 81
rect -264 75 -262 79
rect -728 46 -726 49
rect -692 46 -690 49
rect -684 46 -682 49
rect -648 46 -646 49
rect -640 46 -638 49
rect -597 46 -595 49
rect -515 46 -513 49
rect -479 46 -477 49
rect -471 46 -469 49
rect -435 46 -433 49
rect -427 46 -425 49
rect -384 46 -382 49
rect -151 74 -149 78
rect 22 85 24 88
rect -227 67 -225 74
rect -194 60 -192 74
rect -227 44 -225 47
rect -194 37 -192 40
rect -264 15 -262 35
rect -18 54 -16 74
rect -8 54 -6 74
rect 965 83 967 103
rect 1307 124 1309 131
rect 1302 120 1309 124
rect 1303 109 1305 120
rect 1315 112 1317 131
rect 1345 123 1347 131
rect 1389 123 1391 131
rect 1339 121 1347 123
rect 1383 121 1391 123
rect 1339 109 1341 121
rect 1347 109 1349 118
rect 1383 109 1385 121
rect 1391 109 1393 118
rect 1434 109 1436 131
rect 1002 95 1004 98
rect 22 59 24 73
rect 697 69 699 76
rect 692 65 699 69
rect 693 54 695 65
rect 705 57 707 76
rect 735 68 737 76
rect 779 68 781 76
rect 729 66 737 68
rect 773 66 781 68
rect 729 54 731 66
rect 737 54 739 63
rect 773 54 775 66
rect 781 54 783 63
rect 824 54 826 76
rect 1035 88 1037 91
rect 965 60 967 63
rect 1002 61 1004 75
rect 1078 82 1080 102
rect 1303 96 1305 99
rect 1339 96 1341 99
rect 1347 96 1349 99
rect 1383 96 1385 99
rect 1391 96 1393 99
rect 1434 96 1436 99
rect 1035 61 1037 68
rect 1078 59 1080 62
rect 22 50 24 53
rect -18 39 -16 42
rect -8 39 -6 42
rect 693 41 695 44
rect 729 41 731 44
rect 737 41 739 44
rect 773 41 775 44
rect 781 41 783 44
rect 824 41 826 44
rect -227 27 -225 30
rect -194 20 -192 23
rect -264 -8 -262 -5
rect -227 -7 -225 7
rect -151 14 -149 34
rect 511 32 513 35
rect 521 32 523 35
rect 265 21 267 25
rect -194 -7 -192 0
rect -151 -9 -149 -6
rect 378 20 380 24
rect 551 31 553 34
rect 302 13 304 20
rect 335 6 337 20
rect 302 -10 304 -7
rect 335 -17 337 -14
rect 265 -39 267 -19
rect 511 0 513 20
rect 521 0 523 20
rect 551 5 553 19
rect 551 -4 553 -1
rect 630 -4 632 -1
rect 640 -4 642 -1
rect 511 -15 513 -12
rect 521 -15 523 -12
rect 302 -27 304 -24
rect 335 -34 337 -31
rect 265 -62 267 -59
rect 302 -61 304 -47
rect 378 -40 380 -20
rect 671 -17 673 -14
rect 335 -61 337 -54
rect 516 -42 518 -39
rect 526 -42 528 -39
rect 556 -43 558 -40
rect 378 -63 380 -60
rect 516 -74 518 -54
rect 526 -74 528 -54
rect 630 -49 632 -28
rect 640 -49 642 -28
rect 671 -43 673 -29
rect 671 -52 673 -49
rect 556 -69 558 -55
rect 630 -58 632 -55
rect 640 -58 642 -55
rect 556 -78 558 -75
rect 516 -89 518 -86
rect 526 -89 528 -86
rect 1297 -152 1299 -149
rect 1305 -152 1307 -149
rect 1335 -152 1337 -149
rect 1379 -152 1381 -149
rect 1424 -152 1426 -149
rect 955 -165 957 -161
rect 506 -173 508 -170
rect 516 -173 518 -170
rect 260 -184 262 -180
rect -709 -223 -707 -220
rect -701 -223 -699 -220
rect -671 -223 -669 -220
rect -627 -223 -625 -220
rect -582 -223 -580 -220
rect -496 -223 -494 -220
rect -488 -223 -486 -220
rect -458 -223 -456 -220
rect -414 -223 -412 -220
rect -369 -223 -367 -220
rect 373 -185 375 -181
rect 546 -174 548 -171
rect 297 -192 299 -185
rect 330 -199 332 -185
rect 297 -215 299 -212
rect 330 -222 332 -219
rect -3 -243 -1 -240
rect 7 -243 9 -240
rect -709 -255 -707 -248
rect -714 -259 -707 -255
rect -713 -270 -711 -259
rect -701 -267 -699 -248
rect -671 -256 -669 -248
rect -627 -256 -625 -248
rect -677 -258 -669 -256
rect -633 -258 -625 -256
rect -677 -270 -675 -258
rect -669 -270 -667 -261
rect -633 -270 -631 -258
rect -625 -270 -623 -261
rect -582 -270 -580 -248
rect -496 -255 -494 -248
rect -501 -259 -494 -255
rect -500 -270 -498 -259
rect -488 -267 -486 -248
rect -458 -256 -456 -248
rect -414 -256 -412 -248
rect -464 -258 -456 -256
rect -420 -258 -412 -256
rect -464 -270 -462 -258
rect -456 -270 -454 -261
rect -420 -270 -418 -258
rect -412 -270 -410 -261
rect -369 -270 -367 -248
rect -249 -254 -247 -250
rect -713 -283 -711 -280
rect -677 -283 -675 -280
rect -669 -283 -667 -280
rect -633 -283 -631 -280
rect -625 -283 -623 -280
rect -582 -283 -580 -280
rect -500 -283 -498 -280
rect -464 -283 -462 -280
rect -456 -283 -454 -280
rect -420 -283 -418 -280
rect -412 -283 -410 -280
rect -369 -283 -367 -280
rect -136 -255 -134 -251
rect 37 -244 39 -241
rect 260 -244 262 -224
rect 506 -205 508 -185
rect 516 -205 518 -185
rect 546 -200 548 -186
rect 1068 -166 1070 -162
rect 992 -173 994 -166
rect 1025 -180 1027 -166
rect 992 -196 994 -193
rect 1025 -203 1027 -200
rect 546 -209 548 -206
rect 625 -209 627 -206
rect 635 -209 637 -206
rect 506 -220 508 -217
rect 516 -220 518 -217
rect 297 -232 299 -229
rect -212 -262 -210 -255
rect -179 -269 -177 -255
rect -212 -285 -210 -282
rect -179 -292 -177 -289
rect -249 -314 -247 -294
rect -3 -275 -1 -255
rect 7 -275 9 -255
rect 37 -270 39 -256
rect 330 -239 332 -236
rect 260 -267 262 -264
rect 297 -266 299 -252
rect 373 -245 375 -225
rect 666 -222 668 -219
rect 330 -266 332 -259
rect 511 -247 513 -244
rect 521 -247 523 -244
rect 551 -248 553 -245
rect 373 -268 375 -265
rect 37 -279 39 -276
rect 511 -279 513 -259
rect 521 -279 523 -259
rect 625 -254 627 -233
rect 635 -254 637 -233
rect 955 -225 957 -205
rect 1297 -184 1299 -177
rect 1292 -188 1299 -184
rect 1293 -199 1295 -188
rect 1305 -196 1307 -177
rect 1335 -185 1337 -177
rect 1379 -185 1381 -177
rect 1329 -187 1337 -185
rect 1373 -187 1381 -185
rect 1329 -199 1331 -187
rect 1337 -199 1339 -190
rect 1373 -199 1375 -187
rect 1381 -199 1383 -190
rect 1424 -199 1426 -177
rect 992 -213 994 -210
rect 666 -248 668 -234
rect 1025 -220 1027 -217
rect 955 -248 957 -245
rect 992 -247 994 -233
rect 1068 -226 1070 -206
rect 1293 -212 1295 -209
rect 1329 -212 1331 -209
rect 1337 -212 1339 -209
rect 1373 -212 1375 -209
rect 1381 -212 1383 -209
rect 1424 -212 1426 -209
rect 1025 -247 1027 -240
rect 1068 -249 1070 -246
rect 666 -257 668 -254
rect 551 -274 553 -260
rect 625 -263 627 -260
rect 635 -263 637 -260
rect -3 -290 -1 -287
rect 7 -290 9 -287
rect 551 -283 553 -280
rect 511 -294 513 -291
rect 521 -294 523 -291
rect -212 -302 -210 -299
rect -179 -309 -177 -306
rect -249 -337 -247 -334
rect -212 -336 -210 -322
rect -136 -315 -134 -295
rect -179 -336 -177 -329
rect -136 -338 -134 -335
rect 1321 -411 1323 -408
rect 1329 -411 1331 -408
rect 1359 -411 1361 -408
rect 1403 -411 1405 -408
rect 1448 -411 1450 -408
rect 979 -424 981 -420
rect 555 -427 557 -424
rect 565 -427 567 -424
rect 309 -438 311 -434
rect 422 -439 424 -435
rect 595 -428 597 -425
rect 346 -446 348 -439
rect 379 -453 381 -439
rect 346 -469 348 -466
rect 379 -476 381 -473
rect -685 -490 -683 -487
rect -677 -490 -675 -487
rect -647 -490 -645 -487
rect -603 -490 -601 -487
rect -558 -490 -556 -487
rect -472 -490 -470 -487
rect -464 -490 -462 -487
rect -434 -490 -432 -487
rect -390 -490 -388 -487
rect -345 -490 -343 -487
rect 309 -498 311 -478
rect 555 -459 557 -439
rect 565 -459 567 -439
rect 595 -454 597 -440
rect 595 -463 597 -460
rect 674 -463 676 -460
rect 684 -463 686 -460
rect 555 -474 557 -471
rect 565 -474 567 -471
rect 346 -486 348 -483
rect 21 -510 23 -507
rect 31 -510 33 -507
rect -685 -522 -683 -515
rect -690 -526 -683 -522
rect -689 -537 -687 -526
rect -677 -534 -675 -515
rect -647 -523 -645 -515
rect -603 -523 -601 -515
rect -653 -525 -645 -523
rect -609 -525 -601 -523
rect -653 -537 -651 -525
rect -645 -537 -643 -528
rect -609 -537 -607 -525
rect -601 -537 -599 -528
rect -558 -537 -556 -515
rect -472 -522 -470 -515
rect -477 -526 -470 -522
rect -476 -537 -474 -526
rect -464 -534 -462 -515
rect -434 -523 -432 -515
rect -390 -523 -388 -515
rect -440 -525 -432 -523
rect -396 -525 -388 -523
rect -440 -537 -438 -525
rect -432 -537 -430 -528
rect -396 -537 -394 -525
rect -388 -537 -386 -528
rect -345 -537 -343 -515
rect -225 -521 -223 -517
rect -689 -550 -687 -547
rect -653 -550 -651 -547
rect -645 -550 -643 -547
rect -609 -550 -607 -547
rect -601 -550 -599 -547
rect -558 -550 -556 -547
rect -476 -550 -474 -547
rect -440 -550 -438 -547
rect -432 -550 -430 -547
rect -396 -550 -394 -547
rect -388 -550 -386 -547
rect -345 -550 -343 -547
rect -112 -522 -110 -518
rect 61 -511 63 -508
rect -188 -529 -186 -522
rect -155 -536 -153 -522
rect -188 -552 -186 -549
rect -155 -559 -153 -556
rect -225 -581 -223 -561
rect 21 -542 23 -522
rect 31 -542 33 -522
rect 379 -493 381 -490
rect 309 -521 311 -518
rect 346 -520 348 -506
rect 422 -499 424 -479
rect 1092 -425 1094 -421
rect 1016 -432 1018 -425
rect 1049 -439 1051 -425
rect 1016 -455 1018 -452
rect 1049 -462 1051 -459
rect 715 -476 717 -473
rect 379 -520 381 -513
rect 560 -501 562 -498
rect 570 -501 572 -498
rect 600 -502 602 -499
rect 61 -537 63 -523
rect 422 -522 424 -519
rect 560 -533 562 -513
rect 570 -533 572 -513
rect 674 -508 676 -487
rect 684 -508 686 -487
rect 979 -484 981 -464
rect 1321 -443 1323 -436
rect 1316 -447 1323 -443
rect 1317 -458 1319 -447
rect 1329 -455 1331 -436
rect 1359 -444 1361 -436
rect 1403 -444 1405 -436
rect 1353 -446 1361 -444
rect 1397 -446 1405 -444
rect 1353 -458 1355 -446
rect 1361 -458 1363 -449
rect 1397 -458 1399 -446
rect 1405 -458 1407 -449
rect 1448 -458 1450 -436
rect 1016 -472 1018 -469
rect 715 -502 717 -488
rect 1049 -479 1051 -476
rect 979 -507 981 -504
rect 1016 -506 1018 -492
rect 1092 -485 1094 -465
rect 1317 -471 1319 -468
rect 1353 -471 1355 -468
rect 1361 -471 1363 -468
rect 1397 -471 1399 -468
rect 1405 -471 1407 -468
rect 1448 -471 1450 -468
rect 1049 -506 1051 -499
rect 715 -511 717 -508
rect 1092 -508 1094 -505
rect 600 -528 602 -514
rect 674 -517 676 -514
rect 684 -517 686 -514
rect 61 -546 63 -543
rect 600 -537 602 -534
rect 560 -548 562 -545
rect 570 -548 572 -545
rect 21 -557 23 -554
rect 31 -557 33 -554
rect -188 -569 -186 -566
rect -155 -576 -153 -573
rect -225 -604 -223 -601
rect -188 -603 -186 -589
rect -112 -582 -110 -562
rect -155 -603 -153 -596
rect -112 -605 -110 -602
rect 550 -632 552 -629
rect 560 -632 562 -629
rect 304 -643 306 -639
rect 417 -644 419 -640
rect 590 -633 592 -630
rect 341 -651 343 -644
rect 374 -658 376 -644
rect 341 -674 343 -671
rect 374 -681 376 -678
rect 304 -703 306 -683
rect 550 -664 552 -644
rect 560 -664 562 -644
rect 590 -659 592 -645
rect 590 -668 592 -665
rect 669 -668 671 -665
rect 679 -668 681 -665
rect 550 -679 552 -676
rect 560 -679 562 -676
rect 341 -691 343 -688
rect 374 -698 376 -695
rect 304 -726 306 -723
rect 341 -725 343 -711
rect 417 -704 419 -684
rect 750 -677 752 -674
rect 758 -677 760 -674
rect 788 -677 790 -674
rect 832 -677 834 -674
rect 877 -677 879 -674
rect 710 -681 712 -678
rect 374 -725 376 -718
rect 555 -706 557 -703
rect 565 -706 567 -703
rect 595 -707 597 -704
rect 417 -727 419 -724
rect 555 -738 557 -718
rect 565 -738 567 -718
rect 669 -713 671 -692
rect 679 -713 681 -692
rect 710 -707 712 -693
rect 750 -709 752 -702
rect 745 -713 752 -709
rect 710 -716 712 -713
rect 595 -733 597 -719
rect 669 -722 671 -719
rect 679 -722 681 -719
rect 746 -724 748 -713
rect 758 -721 760 -702
rect 788 -710 790 -702
rect 832 -710 834 -702
rect 782 -712 790 -710
rect 826 -712 834 -710
rect 782 -724 784 -712
rect 790 -724 792 -715
rect 826 -724 828 -712
rect 834 -724 836 -715
rect 877 -724 879 -702
rect 1342 -717 1344 -714
rect 1350 -717 1352 -714
rect 1380 -717 1382 -714
rect 1424 -717 1426 -714
rect 1469 -717 1471 -714
rect 1000 -730 1002 -726
rect 746 -737 748 -734
rect 782 -737 784 -734
rect 790 -737 792 -734
rect 826 -737 828 -734
rect 834 -737 836 -734
rect 877 -737 879 -734
rect 595 -742 597 -739
rect 555 -753 557 -750
rect 565 -753 567 -750
rect 1113 -731 1115 -727
rect 1037 -738 1039 -731
rect 1070 -745 1072 -731
rect 1037 -761 1039 -758
rect 1070 -768 1072 -765
rect 1000 -790 1002 -770
rect 1342 -749 1344 -742
rect 1337 -753 1344 -749
rect 1338 -764 1340 -753
rect 1350 -761 1352 -742
rect 1380 -750 1382 -742
rect 1424 -750 1426 -742
rect 1374 -752 1382 -750
rect 1418 -752 1426 -750
rect 1374 -764 1376 -752
rect 1382 -764 1384 -755
rect 1418 -764 1420 -752
rect 1426 -764 1428 -755
rect 1469 -764 1471 -742
rect 1037 -778 1039 -775
rect -656 -800 -654 -797
rect -648 -800 -646 -797
rect -618 -800 -616 -797
rect -574 -800 -572 -797
rect -529 -800 -527 -797
rect -443 -800 -441 -797
rect -435 -800 -433 -797
rect -405 -800 -403 -797
rect -361 -800 -359 -797
rect -316 -800 -314 -797
rect 1070 -785 1072 -782
rect 1000 -813 1002 -810
rect 1037 -812 1039 -798
rect 1113 -791 1115 -771
rect 1338 -777 1340 -774
rect 1374 -777 1376 -774
rect 1382 -777 1384 -774
rect 1418 -777 1420 -774
rect 1426 -777 1428 -774
rect 1469 -777 1471 -774
rect 1070 -812 1072 -805
rect 1113 -814 1115 -811
rect 50 -820 52 -817
rect 60 -820 62 -817
rect -656 -832 -654 -825
rect -661 -836 -654 -832
rect -660 -847 -658 -836
rect -648 -844 -646 -825
rect -618 -833 -616 -825
rect -574 -833 -572 -825
rect -624 -835 -616 -833
rect -580 -835 -572 -833
rect -624 -847 -622 -835
rect -616 -847 -614 -838
rect -580 -847 -578 -835
rect -572 -847 -570 -838
rect -529 -847 -527 -825
rect -443 -832 -441 -825
rect -448 -836 -441 -832
rect -447 -847 -445 -836
rect -435 -844 -433 -825
rect -405 -833 -403 -825
rect -361 -833 -359 -825
rect -411 -835 -403 -833
rect -367 -835 -359 -833
rect -411 -847 -409 -835
rect -403 -847 -401 -838
rect -367 -847 -365 -835
rect -359 -847 -357 -838
rect -316 -847 -314 -825
rect -196 -831 -194 -827
rect -660 -860 -658 -857
rect -624 -860 -622 -857
rect -616 -860 -614 -857
rect -580 -860 -578 -857
rect -572 -860 -570 -857
rect -529 -860 -527 -857
rect -447 -860 -445 -857
rect -411 -860 -409 -857
rect -403 -860 -401 -857
rect -367 -860 -365 -857
rect -359 -860 -357 -857
rect -316 -860 -314 -857
rect -83 -832 -81 -828
rect 90 -821 92 -818
rect -159 -839 -157 -832
rect -126 -846 -124 -832
rect -159 -862 -157 -859
rect -126 -869 -124 -866
rect -196 -891 -194 -871
rect 50 -852 52 -832
rect 60 -852 62 -832
rect 90 -847 92 -833
rect 90 -856 92 -853
rect 50 -867 52 -864
rect 60 -867 62 -864
rect -159 -879 -157 -876
rect -126 -886 -124 -883
rect -196 -914 -194 -911
rect -159 -913 -157 -899
rect -83 -892 -81 -872
rect -126 -913 -124 -906
rect -83 -915 -81 -912
<< polycontact >>
rect 1001 142 1005 147
rect 1034 142 1038 147
rect -733 70 -729 74
rect -720 62 -716 66
rect -697 62 -692 67
rect -682 62 -677 66
rect -653 62 -648 67
rect -601 67 -597 72
rect -638 62 -633 66
rect -520 70 -516 74
rect -507 62 -503 66
rect -484 62 -479 67
rect -469 62 -464 66
rect -440 62 -435 67
rect -388 67 -384 72
rect -425 62 -420 66
rect -228 74 -224 79
rect -195 74 -191 79
rect -268 18 -264 23
rect -22 63 -18 67
rect -12 57 -8 61
rect 961 86 965 91
rect 1298 120 1302 124
rect 1311 112 1315 116
rect 1334 112 1339 117
rect 1349 112 1354 116
rect 1378 112 1383 117
rect 1430 117 1434 122
rect 1393 112 1398 116
rect 18 62 22 66
rect 688 65 692 69
rect 701 57 705 61
rect 724 57 729 62
rect 739 57 744 61
rect 768 57 773 62
rect 820 62 824 67
rect 783 57 788 61
rect 1074 85 1078 90
rect 1001 56 1005 61
rect 1034 56 1038 61
rect -155 17 -151 22
rect -228 -12 -224 -7
rect -195 -12 -191 -7
rect 301 20 305 25
rect 334 20 338 25
rect 261 -36 265 -31
rect 507 9 511 13
rect 517 3 521 7
rect 547 8 551 12
rect 374 -37 378 -32
rect 301 -66 305 -61
rect 334 -66 338 -61
rect 512 -65 516 -61
rect 522 -71 526 -67
rect 626 -46 630 -42
rect 636 -39 640 -35
rect 667 -40 671 -36
rect 552 -66 556 -62
rect 296 -185 300 -180
rect 329 -185 333 -180
rect 256 -241 260 -236
rect -718 -259 -714 -255
rect -705 -267 -701 -263
rect -682 -267 -677 -262
rect -667 -267 -662 -263
rect -638 -267 -633 -262
rect -586 -262 -582 -257
rect -623 -267 -618 -263
rect -505 -259 -501 -255
rect -492 -267 -488 -263
rect -469 -267 -464 -262
rect -454 -267 -449 -263
rect -425 -267 -420 -262
rect -373 -262 -369 -257
rect -410 -267 -405 -263
rect -213 -255 -209 -250
rect -180 -255 -176 -250
rect 502 -196 506 -192
rect 512 -202 516 -198
rect 542 -197 546 -193
rect 991 -166 995 -161
rect 1024 -166 1028 -161
rect -253 -311 -249 -306
rect -7 -266 -3 -262
rect 3 -272 7 -268
rect 33 -267 37 -263
rect 369 -242 373 -237
rect 951 -222 955 -217
rect 296 -271 300 -266
rect 329 -271 333 -266
rect 507 -270 511 -266
rect 517 -276 521 -272
rect 621 -251 625 -247
rect 631 -244 635 -240
rect 1288 -188 1292 -184
rect 1301 -196 1305 -192
rect 1324 -196 1329 -191
rect 1339 -196 1344 -192
rect 1368 -196 1373 -191
rect 1420 -191 1424 -186
rect 1383 -196 1388 -192
rect 662 -245 666 -241
rect 1064 -223 1068 -218
rect 991 -252 995 -247
rect 1024 -252 1028 -247
rect 547 -271 551 -267
rect -140 -312 -136 -307
rect -213 -341 -209 -336
rect -180 -341 -176 -336
rect 345 -439 349 -434
rect 378 -439 382 -434
rect 305 -495 309 -490
rect 551 -450 555 -446
rect 561 -456 565 -452
rect 591 -451 595 -447
rect -694 -526 -690 -522
rect -681 -534 -677 -530
rect -658 -534 -653 -529
rect -643 -534 -638 -530
rect -614 -534 -609 -529
rect -562 -529 -558 -524
rect -599 -534 -594 -530
rect -481 -526 -477 -522
rect -468 -534 -464 -530
rect -445 -534 -440 -529
rect -430 -534 -425 -530
rect -401 -534 -396 -529
rect -349 -529 -345 -524
rect -386 -534 -381 -530
rect -189 -522 -185 -517
rect -156 -522 -152 -517
rect -229 -578 -225 -573
rect 17 -533 21 -529
rect 27 -539 31 -535
rect 418 -496 422 -491
rect 1015 -425 1019 -420
rect 1048 -425 1052 -420
rect 57 -534 61 -530
rect 345 -525 349 -520
rect 378 -525 382 -520
rect 556 -524 560 -520
rect 566 -530 570 -526
rect 670 -505 674 -501
rect 680 -498 684 -494
rect 975 -481 979 -476
rect 1312 -447 1316 -443
rect 1325 -455 1329 -451
rect 1348 -455 1353 -450
rect 1363 -455 1368 -451
rect 1392 -455 1397 -450
rect 1444 -450 1448 -445
rect 1407 -455 1412 -451
rect 711 -499 715 -495
rect 1088 -482 1092 -477
rect 1015 -511 1019 -506
rect 1048 -511 1052 -506
rect 596 -525 600 -521
rect -116 -579 -112 -574
rect -189 -608 -185 -603
rect -156 -608 -152 -603
rect 340 -644 344 -639
rect 373 -644 377 -639
rect 300 -700 304 -695
rect 546 -655 550 -651
rect 556 -661 560 -657
rect 586 -656 590 -652
rect 413 -701 417 -696
rect 340 -730 344 -725
rect 373 -730 377 -725
rect 551 -729 555 -725
rect 561 -735 565 -731
rect 665 -710 669 -706
rect 675 -703 679 -699
rect 706 -704 710 -700
rect 741 -713 745 -709
rect 591 -730 595 -726
rect 754 -721 758 -717
rect 777 -721 782 -716
rect 792 -721 797 -717
rect 821 -721 826 -716
rect 873 -716 877 -711
rect 836 -721 841 -717
rect 1036 -731 1040 -726
rect 1069 -731 1073 -726
rect 996 -787 1000 -782
rect 1333 -753 1337 -749
rect 1346 -761 1350 -757
rect 1369 -761 1374 -756
rect 1384 -761 1389 -757
rect 1413 -761 1418 -756
rect 1465 -756 1469 -751
rect 1428 -761 1433 -757
rect 1109 -788 1113 -783
rect 1036 -817 1040 -812
rect 1069 -817 1073 -812
rect -665 -836 -661 -832
rect -652 -844 -648 -840
rect -629 -844 -624 -839
rect -614 -844 -609 -840
rect -585 -844 -580 -839
rect -533 -839 -529 -834
rect -570 -844 -565 -840
rect -452 -836 -448 -832
rect -439 -844 -435 -840
rect -416 -844 -411 -839
rect -401 -844 -396 -840
rect -372 -844 -367 -839
rect -320 -839 -316 -834
rect -357 -844 -352 -840
rect -160 -832 -156 -827
rect -127 -832 -123 -827
rect -200 -888 -196 -883
rect 46 -843 50 -839
rect 56 -849 60 -845
rect 86 -844 90 -840
rect -87 -889 -83 -884
rect -160 -918 -156 -913
rect -127 -918 -123 -913
<< metal1 >>
rect 932 179 1165 184
rect 960 143 964 179
rect -735 112 -31 116
rect -729 106 -725 112
rect -691 106 -687 112
rect -647 106 -643 112
rect -602 106 -598 112
rect -516 106 -512 112
rect -478 106 -474 112
rect -434 106 -430 112
rect -389 106 -385 112
rect -297 111 -31 112
rect -679 81 -666 106
rect -635 81 -622 106
rect -466 81 -453 106
rect -422 81 -409 106
rect -740 70 -733 74
rect -713 73 -709 81
rect -713 70 -673 73
rect -723 62 -720 66
rect -713 59 -709 70
rect -701 62 -697 67
rect -677 62 -673 70
rect -669 67 -666 81
rect -625 72 -622 81
rect -625 67 -601 72
rect -594 71 -590 81
rect -669 62 -653 67
rect -633 62 -629 66
rect -669 59 -666 62
rect -625 59 -622 67
rect -594 66 -581 71
rect -594 59 -590 66
rect -527 70 -520 74
rect -500 73 -496 81
rect -500 70 -460 73
rect -510 62 -507 66
rect -500 59 -496 70
rect -488 62 -484 67
rect -464 62 -460 70
rect -456 67 -453 81
rect -412 72 -409 81
rect -412 67 -388 72
rect -381 71 -377 81
rect -269 75 -265 111
rect -456 62 -440 67
rect -420 62 -416 66
rect -456 59 -453 62
rect -412 59 -409 67
rect -381 66 -368 71
rect -381 59 -377 66
rect -721 49 -709 59
rect -677 49 -666 59
rect -633 49 -622 59
rect -508 49 -496 59
rect -464 49 -453 59
rect -420 49 -409 59
rect -733 44 -729 49
rect -697 44 -693 49
rect -653 44 -649 49
rect -602 44 -598 49
rect -520 44 -516 49
rect -484 44 -480 49
rect -440 44 -436 49
rect -389 44 -385 49
rect -734 40 -377 44
rect -381 -45 -377 40
rect -244 43 -239 98
rect -228 79 -224 86
rect -195 79 -191 86
rect -156 74 -152 111
rect -69 91 -63 98
rect -36 95 -31 111
rect 686 107 839 111
rect 692 101 696 107
rect 730 101 734 107
rect 774 101 778 107
rect 819 101 823 107
rect 985 111 990 166
rect 1001 147 1005 154
rect 1034 147 1038 154
rect 1073 142 1077 179
rect 1120 159 1171 165
rect 1296 162 1449 166
rect 1093 154 1171 159
rect 1302 156 1306 162
rect 1340 156 1344 162
rect 1384 156 1388 162
rect 1429 156 1433 162
rect 997 111 1001 115
rect 985 107 1001 111
rect -36 94 14 95
rect -36 92 35 94
rect -136 86 -55 91
rect -232 43 -228 47
rect -244 39 -228 43
rect -278 18 -268 23
rect -261 22 -257 35
rect -232 27 -228 39
rect -261 17 -248 22
rect -261 15 -257 17
rect -224 42 -220 47
rect -224 38 -207 42
rect -224 27 -220 38
rect -211 28 -207 38
rect -199 28 -195 40
rect -211 23 -195 28
rect -269 -44 -265 -5
rect -228 -25 -224 -12
rect -211 -38 -205 23
rect -199 20 -195 23
rect -191 27 -187 40
rect -191 23 -170 27
rect -191 20 -187 23
rect -176 22 -170 23
rect -176 17 -166 22
rect -160 17 -155 22
rect -148 21 -144 34
rect -106 60 -97 73
rect -58 66 -55 86
rect -23 86 -20 92
rect -4 86 -1 92
rect 11 91 35 92
rect 17 85 20 91
rect -14 71 -11 74
rect 742 76 755 101
rect 786 76 799 101
rect 951 86 961 91
rect 968 90 972 103
rect 997 95 1001 107
rect 968 85 981 90
rect 968 83 972 85
rect -14 68 -1 71
rect -58 63 -22 66
rect -4 65 -1 68
rect -4 62 18 65
rect 26 65 29 73
rect 681 65 688 69
rect 708 68 712 76
rect 708 65 748 68
rect 26 62 38 65
rect -106 57 -12 60
rect -148 16 -131 21
rect -148 14 -144 16
rect -195 -25 -191 -12
rect -156 -44 -152 -6
rect -106 -24 -98 57
rect -4 54 -1 62
rect 26 59 29 62
rect 184 57 498 62
rect 698 57 701 61
rect 17 49 20 53
rect 7 46 35 49
rect -23 36 -20 42
rect 7 36 11 46
rect -88 33 11 36
rect -88 -44 -77 33
rect -297 -45 -77 -44
rect -381 -52 -77 -45
rect 184 -143 190 57
rect 260 21 264 57
rect 285 -11 290 44
rect 301 25 305 32
rect 334 25 338 32
rect 373 20 377 57
rect 493 41 498 57
rect 708 54 712 65
rect 720 57 724 62
rect 744 57 748 65
rect 752 62 755 76
rect 796 67 799 76
rect 796 62 820 67
rect 827 66 831 76
rect 752 57 768 62
rect 788 57 792 61
rect 752 54 755 57
rect 796 54 799 62
rect 827 61 840 66
rect 1005 110 1009 115
rect 1005 106 1022 110
rect 1005 95 1009 106
rect 1018 96 1022 106
rect 1030 96 1034 108
rect 1018 91 1034 96
rect 827 54 831 61
rect 700 44 712 54
rect 744 44 755 54
rect 788 44 799 54
rect 493 40 543 41
rect 493 38 619 40
rect 688 39 692 44
rect 724 39 728 44
rect 768 39 772 44
rect 819 39 823 44
rect 393 32 474 37
rect 297 -11 301 -7
rect 285 -15 301 -11
rect 251 -36 261 -31
rect 268 -32 272 -19
rect 297 -27 301 -15
rect 268 -37 281 -32
rect 268 -39 272 -37
rect 305 -12 309 -7
rect 305 -16 322 -12
rect 305 -27 309 -16
rect 318 -26 322 -16
rect 330 -26 334 -14
rect 318 -31 334 -26
rect 226 -98 237 -97
rect 260 -98 264 -59
rect 301 -79 305 -66
rect 318 -90 324 -31
rect 330 -34 334 -31
rect 338 -27 342 -14
rect 471 12 474 32
rect 493 32 498 38
rect 506 32 509 38
rect 525 32 528 38
rect 540 37 619 38
rect 546 31 549 37
rect 515 17 518 20
rect 515 14 528 17
rect 471 9 507 12
rect 525 11 528 14
rect 525 8 547 11
rect 555 11 558 19
rect 555 8 582 11
rect 338 -31 359 -27
rect 338 -34 342 -31
rect 353 -32 359 -31
rect 353 -37 363 -32
rect 369 -37 374 -32
rect 381 -33 385 -20
rect 423 3 517 6
rect 381 -38 398 -33
rect 381 -40 385 -38
rect 334 -79 338 -66
rect 373 -98 377 -60
rect 423 -78 431 3
rect 525 0 528 8
rect 555 5 558 8
rect 546 -5 549 -1
rect 536 -8 564 -5
rect 506 -18 509 -12
rect 536 -18 540 -8
rect 441 -21 540 -18
rect 441 -98 452 -21
rect 498 -34 548 -33
rect 498 -36 569 -34
rect 511 -42 514 -36
rect 530 -42 533 -36
rect 545 -37 569 -36
rect 579 -36 582 8
rect 615 5 619 37
rect 687 35 831 39
rect 960 24 964 63
rect 1001 43 1005 56
rect 1018 33 1024 91
rect 1030 88 1034 91
rect 1038 95 1042 108
rect 1352 131 1365 156
rect 1396 131 1409 156
rect 1281 120 1298 124
rect 1318 123 1322 131
rect 1318 120 1358 123
rect 1308 112 1311 116
rect 1318 109 1322 120
rect 1330 112 1334 117
rect 1354 112 1358 120
rect 1362 117 1365 131
rect 1406 122 1409 131
rect 1406 117 1430 122
rect 1437 121 1441 131
rect 1362 112 1378 117
rect 1398 112 1402 116
rect 1362 109 1365 112
rect 1406 109 1409 117
rect 1437 116 1450 121
rect 1437 109 1441 116
rect 1038 91 1059 95
rect 1038 88 1042 91
rect 1053 90 1059 91
rect 1053 85 1063 90
rect 1069 85 1074 90
rect 1081 89 1085 102
rect 1310 99 1322 109
rect 1354 99 1365 109
rect 1398 99 1409 109
rect 1298 94 1302 99
rect 1334 94 1338 99
rect 1378 94 1382 99
rect 1429 94 1433 99
rect 1297 90 1441 94
rect 1081 84 1098 89
rect 1081 82 1085 84
rect 1123 81 1141 87
rect 1034 43 1038 56
rect 1073 24 1077 62
rect 1123 44 1131 81
rect 932 16 1141 24
rect 615 2 661 5
rect 625 -4 628 2
rect 658 -8 661 2
rect 658 -11 684 -8
rect 551 -43 554 -37
rect 579 -39 636 -36
rect 644 -37 647 -28
rect 666 -17 669 -11
rect 644 -40 667 -37
rect 675 -37 678 -29
rect 675 -40 695 -37
rect 520 -57 523 -54
rect 520 -60 533 -57
rect 503 -65 512 -62
rect 530 -63 533 -60
rect 530 -66 552 -63
rect 560 -63 563 -55
rect 602 -45 626 -42
rect 602 -63 606 -45
rect 644 -43 647 -40
rect 675 -43 678 -40
rect 635 -46 647 -43
rect 635 -49 638 -46
rect 666 -53 669 -49
rect 625 -61 628 -55
rect 644 -61 647 -55
rect 656 -56 684 -53
rect 656 -61 660 -56
rect 560 -66 606 -63
rect 616 -64 660 -61
rect 482 -71 522 -68
rect 482 -90 488 -71
rect 530 -74 533 -66
rect 560 -69 563 -66
rect 551 -79 554 -75
rect 616 -79 619 -64
rect 541 -82 619 -79
rect 511 -92 514 -86
rect 541 -92 545 -82
rect 690 -86 695 -40
rect 500 -95 545 -92
rect 226 -101 452 -98
rect 500 -101 503 -95
rect 226 -106 503 -101
rect 922 -129 1155 -124
rect 184 -148 493 -143
rect -720 -217 -16 -213
rect -714 -223 -710 -217
rect -676 -223 -672 -217
rect -632 -223 -628 -217
rect -587 -223 -583 -217
rect -501 -223 -497 -217
rect -463 -223 -459 -217
rect -419 -223 -415 -217
rect -374 -223 -370 -217
rect -282 -218 -16 -217
rect -664 -248 -651 -223
rect -620 -248 -607 -223
rect -451 -248 -438 -223
rect -407 -248 -394 -223
rect -725 -259 -718 -255
rect -698 -256 -694 -248
rect -698 -259 -658 -256
rect -708 -267 -705 -263
rect -698 -270 -694 -259
rect -686 -267 -682 -262
rect -662 -267 -658 -259
rect -654 -262 -651 -248
rect -610 -257 -607 -248
rect -610 -262 -586 -257
rect -579 -258 -575 -248
rect -654 -267 -638 -262
rect -618 -267 -614 -263
rect -654 -270 -651 -267
rect -610 -270 -607 -262
rect -579 -263 -566 -258
rect -579 -270 -575 -263
rect -512 -259 -505 -255
rect -485 -256 -481 -248
rect -485 -259 -445 -256
rect -495 -267 -492 -263
rect -485 -270 -481 -259
rect -473 -267 -469 -262
rect -449 -267 -445 -259
rect -441 -262 -438 -248
rect -397 -257 -394 -248
rect -397 -262 -373 -257
rect -366 -258 -362 -248
rect -254 -254 -250 -218
rect -441 -267 -425 -262
rect -405 -267 -401 -263
rect -441 -270 -438 -267
rect -397 -270 -394 -262
rect -366 -263 -353 -258
rect -366 -270 -362 -263
rect -706 -280 -694 -270
rect -662 -280 -651 -270
rect -618 -280 -607 -270
rect -493 -280 -481 -270
rect -449 -280 -438 -270
rect -405 -280 -394 -270
rect -718 -285 -714 -280
rect -682 -285 -678 -280
rect -638 -285 -634 -280
rect -587 -285 -583 -280
rect -505 -285 -501 -280
rect -469 -285 -465 -280
rect -425 -285 -421 -280
rect -374 -285 -370 -280
rect -719 -289 -362 -285
rect -366 -374 -362 -289
rect -229 -286 -224 -231
rect -213 -250 -209 -243
rect -180 -250 -176 -243
rect -141 -255 -137 -218
rect -54 -238 -48 -231
rect -21 -234 -16 -218
rect -21 -235 29 -234
rect -21 -237 50 -235
rect -121 -243 -40 -238
rect -217 -286 -213 -282
rect -229 -290 -213 -286
rect -263 -311 -253 -306
rect -246 -307 -242 -294
rect -217 -302 -213 -290
rect -246 -312 -233 -307
rect -246 -314 -242 -312
rect -209 -287 -205 -282
rect -209 -291 -192 -287
rect -209 -302 -205 -291
rect -196 -301 -192 -291
rect -184 -301 -180 -289
rect -196 -306 -180 -301
rect -254 -373 -250 -334
rect -213 -354 -209 -341
rect -196 -367 -190 -306
rect -184 -309 -180 -306
rect -176 -302 -172 -289
rect -176 -306 -155 -302
rect -176 -309 -172 -306
rect -161 -307 -155 -306
rect -161 -312 -151 -307
rect -145 -312 -140 -307
rect -133 -308 -129 -295
rect -91 -269 -82 -256
rect -43 -263 -40 -243
rect -8 -243 -5 -237
rect 11 -243 14 -237
rect 26 -238 50 -237
rect 32 -244 35 -238
rect 1 -258 4 -255
rect 1 -261 14 -258
rect -43 -266 -7 -263
rect 11 -264 14 -261
rect 11 -267 33 -264
rect 41 -264 44 -256
rect 41 -267 53 -264
rect -91 -272 3 -269
rect -133 -313 -116 -308
rect -133 -315 -129 -313
rect -180 -354 -176 -341
rect -141 -373 -137 -335
rect -91 -353 -83 -272
rect 11 -275 14 -267
rect 41 -270 44 -267
rect 32 -280 35 -276
rect 22 -283 50 -280
rect -8 -293 -5 -287
rect 22 -293 26 -283
rect -73 -296 26 -293
rect -73 -373 -62 -296
rect -282 -374 -62 -373
rect -366 -381 -62 -374
rect 184 -397 190 -148
rect 255 -184 259 -148
rect 280 -216 285 -161
rect 296 -180 300 -173
rect 329 -180 333 -173
rect 368 -185 372 -148
rect 488 -164 493 -148
rect 488 -165 538 -164
rect 950 -165 954 -129
rect 488 -167 614 -165
rect 388 -173 469 -168
rect 292 -216 296 -212
rect 280 -220 296 -216
rect 246 -241 256 -236
rect 263 -237 267 -224
rect 292 -232 296 -220
rect 263 -242 276 -237
rect 263 -244 267 -242
rect 215 -303 220 -251
rect 300 -217 304 -212
rect 300 -221 317 -217
rect 300 -232 304 -221
rect 313 -231 317 -221
rect 325 -231 329 -219
rect 313 -236 329 -231
rect 255 -303 259 -264
rect 296 -284 300 -271
rect 313 -295 319 -236
rect 325 -239 329 -236
rect 333 -232 337 -219
rect 466 -193 469 -173
rect 488 -173 493 -167
rect 501 -173 504 -167
rect 520 -173 523 -167
rect 535 -168 614 -167
rect 541 -174 544 -168
rect 510 -188 513 -185
rect 510 -191 523 -188
rect 466 -196 502 -193
rect 520 -194 523 -191
rect 520 -197 542 -194
rect 550 -194 553 -186
rect 550 -197 577 -194
rect 333 -236 354 -232
rect 333 -239 337 -236
rect 348 -237 354 -236
rect 348 -242 358 -237
rect 364 -242 369 -237
rect 376 -238 380 -225
rect 418 -202 512 -199
rect 376 -243 393 -238
rect 376 -245 380 -243
rect 329 -284 333 -271
rect 368 -303 372 -265
rect 418 -283 426 -202
rect 520 -205 523 -197
rect 550 -200 553 -197
rect 541 -210 544 -206
rect 531 -213 559 -210
rect 501 -223 504 -217
rect 531 -223 535 -213
rect 436 -226 535 -223
rect 436 -303 447 -226
rect 493 -239 543 -238
rect 493 -241 564 -239
rect 506 -247 509 -241
rect 525 -247 528 -241
rect 540 -242 564 -241
rect 574 -241 577 -197
rect 610 -200 614 -168
rect 610 -203 656 -200
rect 620 -209 623 -203
rect 653 -213 656 -203
rect 975 -197 980 -142
rect 991 -161 995 -154
rect 1024 -161 1028 -154
rect 1063 -166 1067 -129
rect 1110 -149 1161 -143
rect 1286 -146 1439 -142
rect 1083 -154 1161 -149
rect 1292 -152 1296 -146
rect 1330 -152 1334 -146
rect 1374 -152 1378 -146
rect 1419 -152 1423 -146
rect 987 -197 991 -193
rect 975 -201 991 -197
rect 653 -216 679 -213
rect 546 -248 549 -242
rect 574 -244 631 -241
rect 639 -242 642 -233
rect 661 -222 664 -216
rect 941 -222 951 -217
rect 958 -218 962 -205
rect 987 -213 991 -201
rect 958 -223 971 -218
rect 958 -225 962 -223
rect 639 -245 662 -242
rect 670 -242 673 -234
rect 670 -245 693 -242
rect 515 -262 518 -259
rect 515 -265 528 -262
rect 483 -270 507 -267
rect 525 -268 528 -265
rect 525 -271 547 -268
rect 555 -268 558 -260
rect 597 -250 621 -247
rect 597 -268 601 -250
rect 639 -248 642 -245
rect 670 -248 673 -245
rect 630 -251 642 -248
rect 630 -254 633 -251
rect 661 -258 664 -254
rect 620 -266 623 -260
rect 639 -266 642 -260
rect 651 -261 679 -258
rect 651 -266 655 -261
rect 555 -271 601 -268
rect 611 -269 655 -266
rect 477 -276 517 -273
rect 477 -295 483 -276
rect 525 -279 528 -271
rect 555 -274 558 -271
rect 546 -284 549 -280
rect 611 -284 614 -269
rect 536 -287 614 -284
rect 506 -297 509 -291
rect 536 -297 540 -287
rect 688 -291 693 -245
rect 995 -198 999 -193
rect 995 -202 1012 -198
rect 995 -213 999 -202
rect 1008 -212 1012 -202
rect 1020 -212 1024 -200
rect 1008 -217 1024 -212
rect 950 -284 954 -245
rect 991 -265 995 -252
rect 1008 -275 1014 -217
rect 1020 -220 1024 -217
rect 1028 -213 1032 -200
rect 1342 -177 1355 -152
rect 1386 -177 1399 -152
rect 1271 -188 1288 -184
rect 1308 -185 1312 -177
rect 1308 -188 1348 -185
rect 1298 -196 1301 -192
rect 1308 -199 1312 -188
rect 1320 -196 1324 -191
rect 1344 -196 1348 -188
rect 1352 -191 1355 -177
rect 1396 -186 1399 -177
rect 1396 -191 1420 -186
rect 1427 -187 1431 -177
rect 1352 -196 1368 -191
rect 1388 -196 1392 -192
rect 1352 -199 1355 -196
rect 1396 -199 1399 -191
rect 1427 -192 1440 -187
rect 1427 -199 1431 -192
rect 1028 -217 1049 -213
rect 1028 -220 1032 -217
rect 1043 -218 1049 -217
rect 1043 -223 1053 -218
rect 1059 -223 1064 -218
rect 1071 -219 1075 -206
rect 1300 -209 1312 -199
rect 1344 -209 1355 -199
rect 1388 -209 1399 -199
rect 1288 -214 1292 -209
rect 1324 -214 1328 -209
rect 1368 -214 1372 -209
rect 1419 -214 1423 -209
rect 1287 -218 1431 -214
rect 1071 -224 1088 -219
rect 1071 -226 1075 -224
rect 1113 -227 1131 -221
rect 1024 -265 1028 -252
rect 1063 -284 1067 -246
rect 1113 -264 1121 -227
rect 922 -292 1131 -284
rect 495 -300 540 -297
rect 215 -306 447 -303
rect 495 -306 498 -300
rect 215 -311 498 -306
rect 946 -388 1179 -383
rect 184 -402 542 -397
rect 184 -403 234 -402
rect -696 -484 8 -480
rect -690 -490 -686 -484
rect -652 -490 -648 -484
rect -608 -490 -604 -484
rect -563 -490 -559 -484
rect -477 -490 -473 -484
rect -439 -490 -435 -484
rect -395 -490 -391 -484
rect -350 -490 -346 -484
rect -258 -485 8 -484
rect -640 -515 -627 -490
rect -596 -515 -583 -490
rect -427 -515 -414 -490
rect -383 -515 -370 -490
rect -701 -526 -694 -522
rect -674 -523 -670 -515
rect -674 -526 -634 -523
rect -684 -534 -681 -530
rect -674 -537 -670 -526
rect -662 -534 -658 -529
rect -638 -534 -634 -526
rect -630 -529 -627 -515
rect -586 -524 -583 -515
rect -586 -529 -562 -524
rect -555 -525 -551 -515
rect -630 -534 -614 -529
rect -594 -534 -590 -530
rect -630 -537 -627 -534
rect -586 -537 -583 -529
rect -555 -530 -542 -525
rect -555 -537 -551 -530
rect -488 -526 -481 -522
rect -461 -523 -457 -515
rect -461 -526 -421 -523
rect -471 -534 -468 -530
rect -461 -537 -457 -526
rect -449 -534 -445 -529
rect -425 -534 -421 -526
rect -417 -529 -414 -515
rect -373 -524 -370 -515
rect -373 -529 -349 -524
rect -342 -525 -338 -515
rect -230 -521 -226 -485
rect -417 -534 -401 -529
rect -381 -534 -377 -530
rect -417 -537 -414 -534
rect -373 -537 -370 -529
rect -342 -530 -329 -525
rect -342 -537 -338 -530
rect -682 -547 -670 -537
rect -638 -547 -627 -537
rect -594 -547 -583 -537
rect -469 -547 -457 -537
rect -425 -547 -414 -537
rect -381 -547 -370 -537
rect -694 -552 -690 -547
rect -658 -552 -654 -547
rect -614 -552 -610 -547
rect -563 -552 -559 -547
rect -481 -552 -477 -547
rect -445 -552 -441 -547
rect -401 -552 -397 -547
rect -350 -552 -346 -547
rect -695 -556 -338 -552
rect -342 -641 -338 -556
rect -205 -553 -200 -498
rect -189 -517 -185 -510
rect -156 -517 -152 -510
rect -117 -522 -113 -485
rect -30 -505 -24 -498
rect 3 -501 8 -485
rect 3 -502 53 -501
rect 3 -504 74 -502
rect -97 -510 -16 -505
rect -193 -553 -189 -549
rect -205 -557 -189 -553
rect -239 -578 -229 -573
rect -222 -574 -218 -561
rect -193 -569 -189 -557
rect -222 -579 -209 -574
rect -222 -581 -218 -579
rect -185 -554 -181 -549
rect -185 -558 -168 -554
rect -185 -569 -181 -558
rect -172 -568 -168 -558
rect -160 -568 -156 -556
rect -172 -573 -156 -568
rect -230 -640 -226 -601
rect -189 -621 -185 -608
rect -172 -634 -166 -573
rect -160 -576 -156 -573
rect -152 -569 -148 -556
rect -152 -573 -131 -569
rect -152 -576 -148 -573
rect -137 -574 -131 -573
rect -137 -579 -127 -574
rect -121 -579 -116 -574
rect -109 -575 -105 -562
rect -67 -536 -58 -523
rect -19 -530 -16 -510
rect 16 -510 19 -504
rect 35 -510 38 -504
rect 50 -505 74 -504
rect 56 -511 59 -505
rect 25 -525 28 -522
rect 25 -528 38 -525
rect -19 -533 17 -530
rect 35 -531 38 -528
rect 35 -534 57 -531
rect 65 -531 68 -523
rect 65 -534 77 -531
rect -67 -539 27 -536
rect -109 -580 -92 -575
rect -109 -582 -105 -580
rect -156 -621 -152 -608
rect -117 -640 -113 -602
rect -67 -620 -59 -539
rect 35 -542 38 -534
rect 65 -537 68 -534
rect 56 -547 59 -543
rect 46 -550 74 -547
rect 16 -560 19 -554
rect 46 -560 50 -550
rect -49 -563 50 -560
rect -49 -640 -38 -563
rect 228 -602 234 -403
rect 304 -438 308 -402
rect 329 -470 334 -415
rect 345 -434 349 -427
rect 378 -434 382 -427
rect 417 -439 421 -402
rect 537 -418 542 -402
rect 537 -419 587 -418
rect 537 -421 663 -419
rect 437 -427 518 -422
rect 341 -470 345 -466
rect 329 -474 345 -470
rect 295 -495 305 -490
rect 312 -491 316 -478
rect 341 -486 345 -474
rect 312 -496 325 -491
rect 312 -498 316 -496
rect 255 -556 263 -509
rect 349 -471 353 -466
rect 349 -475 366 -471
rect 349 -486 353 -475
rect 362 -485 366 -475
rect 374 -485 378 -473
rect 362 -490 378 -485
rect 270 -557 281 -556
rect 304 -557 308 -518
rect 345 -538 349 -525
rect 362 -549 368 -490
rect 374 -493 378 -490
rect 382 -486 386 -473
rect 515 -447 518 -427
rect 537 -427 542 -421
rect 550 -427 553 -421
rect 569 -427 572 -421
rect 584 -422 663 -421
rect 590 -428 593 -422
rect 559 -442 562 -439
rect 559 -445 572 -442
rect 515 -450 551 -447
rect 569 -448 572 -445
rect 569 -451 591 -448
rect 599 -448 602 -440
rect 599 -451 626 -448
rect 382 -490 403 -486
rect 382 -493 386 -490
rect 397 -491 403 -490
rect 397 -496 407 -491
rect 413 -496 418 -491
rect 425 -492 429 -479
rect 467 -456 561 -453
rect 425 -497 442 -492
rect 425 -499 429 -497
rect 378 -538 382 -525
rect 417 -557 421 -519
rect 467 -537 475 -456
rect 569 -459 572 -451
rect 599 -454 602 -451
rect 590 -464 593 -460
rect 580 -467 608 -464
rect 550 -477 553 -471
rect 580 -477 584 -467
rect 485 -480 584 -477
rect 485 -557 496 -480
rect 542 -493 592 -492
rect 542 -495 613 -493
rect 518 -521 525 -509
rect 555 -501 558 -495
rect 574 -501 577 -495
rect 589 -496 613 -495
rect 623 -495 626 -451
rect 659 -454 663 -422
rect 974 -424 978 -388
rect 659 -457 705 -454
rect 669 -463 672 -457
rect 702 -467 705 -457
rect 999 -456 1004 -401
rect 1015 -420 1019 -413
rect 1048 -420 1052 -413
rect 1087 -425 1091 -388
rect 1134 -408 1185 -402
rect 1310 -405 1463 -401
rect 1107 -413 1185 -408
rect 1316 -411 1320 -405
rect 1354 -411 1358 -405
rect 1398 -411 1402 -405
rect 1443 -411 1447 -405
rect 1011 -456 1015 -452
rect 999 -460 1015 -456
rect 702 -470 728 -467
rect 595 -502 598 -496
rect 623 -498 680 -495
rect 688 -496 691 -487
rect 710 -476 713 -470
rect 965 -481 975 -476
rect 982 -477 986 -464
rect 1011 -472 1015 -460
rect 982 -482 995 -477
rect 982 -484 986 -482
rect 688 -499 711 -496
rect 719 -496 722 -488
rect 719 -499 739 -496
rect 564 -516 567 -513
rect 564 -519 577 -516
rect 518 -524 556 -521
rect 574 -522 577 -519
rect 574 -525 596 -522
rect 604 -522 607 -514
rect 646 -504 670 -501
rect 646 -522 650 -504
rect 688 -502 691 -499
rect 719 -502 722 -499
rect 679 -505 691 -502
rect 679 -508 682 -505
rect 710 -512 713 -508
rect 669 -520 672 -514
rect 688 -520 691 -514
rect 700 -515 728 -512
rect 700 -520 704 -515
rect 604 -525 650 -522
rect 660 -523 704 -520
rect 526 -530 566 -527
rect 526 -549 532 -530
rect 574 -533 577 -525
rect 604 -528 607 -525
rect 595 -538 598 -534
rect 660 -538 663 -523
rect 585 -541 663 -538
rect 555 -551 558 -545
rect 585 -551 589 -541
rect 734 -545 739 -499
rect 1019 -457 1023 -452
rect 1019 -461 1036 -457
rect 1019 -472 1023 -461
rect 1032 -471 1036 -461
rect 1044 -471 1048 -459
rect 1032 -476 1048 -471
rect 974 -543 978 -504
rect 1015 -524 1019 -511
rect 1032 -534 1038 -476
rect 1044 -479 1048 -476
rect 1052 -472 1056 -459
rect 1366 -436 1379 -411
rect 1410 -436 1423 -411
rect 1295 -447 1312 -443
rect 1332 -444 1336 -436
rect 1332 -447 1372 -444
rect 1322 -455 1325 -451
rect 1332 -458 1336 -447
rect 1344 -455 1348 -450
rect 1368 -455 1372 -447
rect 1376 -450 1379 -436
rect 1420 -445 1423 -436
rect 1420 -450 1444 -445
rect 1451 -446 1455 -436
rect 1376 -455 1392 -450
rect 1412 -455 1416 -451
rect 1376 -458 1379 -455
rect 1420 -458 1423 -450
rect 1451 -451 1464 -446
rect 1451 -458 1455 -451
rect 1052 -476 1073 -472
rect 1052 -479 1056 -476
rect 1067 -477 1073 -476
rect 1067 -482 1077 -477
rect 1083 -482 1088 -477
rect 1095 -478 1099 -465
rect 1324 -468 1336 -458
rect 1368 -468 1379 -458
rect 1412 -468 1423 -458
rect 1312 -473 1316 -468
rect 1348 -473 1352 -468
rect 1392 -473 1396 -468
rect 1443 -473 1447 -468
rect 1311 -477 1455 -473
rect 1095 -483 1112 -478
rect 1095 -485 1099 -483
rect 1137 -486 1155 -480
rect 1048 -524 1052 -511
rect 1087 -543 1091 -505
rect 1137 -523 1145 -486
rect 946 -551 1155 -543
rect 544 -554 589 -551
rect 270 -560 496 -557
rect 544 -560 547 -554
rect 270 -565 547 -560
rect 228 -607 537 -602
rect -258 -641 -38 -640
rect -342 -648 -38 -641
rect 299 -643 303 -607
rect 324 -675 329 -620
rect 340 -639 344 -632
rect 373 -639 377 -632
rect 412 -644 416 -607
rect 532 -623 537 -607
rect 532 -624 582 -623
rect 532 -626 658 -624
rect 432 -632 513 -627
rect 336 -675 340 -671
rect 324 -679 340 -675
rect 290 -700 300 -695
rect 307 -696 311 -683
rect 336 -691 340 -679
rect 307 -701 320 -696
rect 307 -703 311 -701
rect 259 -762 264 -710
rect 344 -676 348 -671
rect 344 -680 361 -676
rect 344 -691 348 -680
rect 357 -690 361 -680
rect 369 -690 373 -678
rect 357 -695 373 -690
rect 299 -762 303 -723
rect 340 -743 344 -730
rect 357 -754 363 -695
rect 369 -698 373 -695
rect 377 -691 381 -678
rect 510 -652 513 -632
rect 532 -632 537 -626
rect 545 -632 548 -626
rect 564 -632 567 -626
rect 579 -627 658 -626
rect 585 -633 588 -627
rect 554 -647 557 -644
rect 554 -650 567 -647
rect 510 -655 546 -652
rect 564 -653 567 -650
rect 564 -656 586 -653
rect 594 -653 597 -645
rect 594 -656 621 -653
rect 377 -695 398 -691
rect 377 -698 381 -695
rect 392 -696 398 -695
rect 392 -701 402 -696
rect 408 -701 413 -696
rect 420 -697 424 -684
rect 462 -661 556 -658
rect 420 -702 437 -697
rect 420 -704 424 -702
rect 373 -743 377 -730
rect 412 -762 416 -724
rect 462 -742 470 -661
rect 564 -664 567 -656
rect 594 -659 597 -656
rect 585 -669 588 -665
rect 575 -672 603 -669
rect 545 -682 548 -676
rect 575 -682 579 -672
rect 480 -685 579 -682
rect 480 -762 491 -685
rect 537 -698 587 -697
rect 537 -700 608 -698
rect 550 -706 553 -700
rect 569 -706 572 -700
rect 584 -701 608 -700
rect 618 -700 621 -656
rect 654 -659 658 -627
rect 654 -662 700 -659
rect 664 -668 667 -662
rect 697 -672 700 -662
rect 739 -671 892 -667
rect 697 -675 723 -672
rect 590 -707 593 -701
rect 618 -703 675 -700
rect 683 -701 686 -692
rect 705 -681 708 -675
rect 745 -677 749 -671
rect 783 -677 787 -671
rect 827 -677 831 -671
rect 872 -677 876 -671
rect 683 -704 706 -701
rect 714 -701 717 -693
rect 714 -704 730 -701
rect 795 -702 808 -677
rect 839 -702 852 -677
rect 967 -694 1200 -689
rect 559 -721 562 -718
rect 559 -724 572 -721
rect 527 -729 551 -726
rect 569 -727 572 -724
rect 569 -730 591 -727
rect 599 -727 602 -719
rect 641 -709 665 -706
rect 641 -727 645 -709
rect 683 -707 686 -704
rect 714 -707 717 -704
rect 674 -710 686 -707
rect 674 -713 677 -710
rect 725 -709 730 -704
rect 725 -713 741 -709
rect 761 -710 765 -702
rect 761 -713 801 -710
rect 705 -717 708 -713
rect 664 -725 667 -719
rect 683 -725 686 -719
rect 695 -720 723 -717
rect 695 -725 699 -720
rect 751 -721 754 -717
rect 761 -724 765 -713
rect 773 -721 777 -716
rect 797 -721 801 -713
rect 805 -716 808 -702
rect 849 -711 852 -702
rect 849 -716 873 -711
rect 880 -712 884 -702
rect 805 -721 821 -716
rect 841 -721 845 -717
rect 805 -724 808 -721
rect 849 -724 852 -716
rect 880 -717 893 -712
rect 880 -724 884 -717
rect 599 -730 645 -727
rect 655 -728 699 -725
rect 521 -735 561 -732
rect 521 -754 527 -735
rect 569 -738 572 -730
rect 599 -733 602 -730
rect 590 -743 593 -739
rect 655 -743 658 -728
rect 753 -734 765 -724
rect 797 -734 808 -724
rect 841 -734 852 -724
rect 995 -730 999 -694
rect 741 -739 745 -734
rect 777 -739 781 -734
rect 821 -739 825 -734
rect 872 -739 876 -734
rect 740 -743 884 -739
rect 580 -746 658 -743
rect 550 -756 553 -750
rect 580 -756 584 -746
rect 539 -759 584 -756
rect 259 -765 491 -762
rect 539 -765 542 -759
rect 259 -770 542 -765
rect 1020 -762 1025 -707
rect 1036 -726 1040 -719
rect 1069 -726 1073 -719
rect 1108 -731 1112 -694
rect 1155 -714 1206 -708
rect 1331 -711 1484 -707
rect 1128 -719 1206 -714
rect 1337 -717 1341 -711
rect 1375 -717 1379 -711
rect 1419 -717 1423 -711
rect 1464 -717 1468 -711
rect 1032 -762 1036 -758
rect 1020 -766 1036 -762
rect 986 -787 996 -782
rect 1003 -783 1007 -770
rect 1032 -778 1036 -766
rect 1003 -788 1016 -783
rect 1003 -790 1007 -788
rect -667 -794 37 -790
rect -661 -800 -657 -794
rect -623 -800 -619 -794
rect -579 -800 -575 -794
rect -534 -800 -530 -794
rect -448 -800 -444 -794
rect -410 -800 -406 -794
rect -366 -800 -362 -794
rect -321 -800 -317 -794
rect -229 -795 37 -794
rect -611 -825 -598 -800
rect -567 -825 -554 -800
rect -398 -825 -385 -800
rect -354 -825 -341 -800
rect -672 -836 -665 -832
rect -645 -833 -641 -825
rect -645 -836 -605 -833
rect -655 -844 -652 -840
rect -645 -847 -641 -836
rect -633 -844 -629 -839
rect -609 -844 -605 -836
rect -601 -839 -598 -825
rect -557 -834 -554 -825
rect -557 -839 -533 -834
rect -526 -835 -522 -825
rect -601 -844 -585 -839
rect -565 -844 -561 -840
rect -601 -847 -598 -844
rect -557 -847 -554 -839
rect -526 -840 -513 -835
rect -526 -847 -522 -840
rect -459 -836 -452 -832
rect -432 -833 -428 -825
rect -432 -836 -392 -833
rect -442 -844 -439 -840
rect -432 -847 -428 -836
rect -420 -844 -416 -839
rect -396 -844 -392 -836
rect -388 -839 -385 -825
rect -344 -834 -341 -825
rect -344 -839 -320 -834
rect -313 -835 -309 -825
rect -201 -831 -197 -795
rect -388 -844 -372 -839
rect -352 -844 -348 -840
rect -388 -847 -385 -844
rect -344 -847 -341 -839
rect -313 -840 -300 -835
rect -313 -847 -309 -840
rect -653 -857 -641 -847
rect -609 -857 -598 -847
rect -565 -857 -554 -847
rect -440 -857 -428 -847
rect -396 -857 -385 -847
rect -352 -857 -341 -847
rect -665 -862 -661 -857
rect -629 -862 -625 -857
rect -585 -862 -581 -857
rect -534 -862 -530 -857
rect -452 -862 -448 -857
rect -416 -862 -412 -857
rect -372 -862 -368 -857
rect -321 -862 -317 -857
rect -666 -866 -309 -862
rect -313 -951 -309 -866
rect -176 -863 -171 -808
rect -160 -827 -156 -820
rect -127 -827 -123 -820
rect -88 -832 -84 -795
rect -1 -815 5 -808
rect 32 -811 37 -795
rect 1040 -763 1044 -758
rect 1040 -767 1057 -763
rect 1040 -778 1044 -767
rect 1053 -777 1057 -767
rect 1065 -777 1069 -765
rect 1053 -782 1069 -777
rect 32 -812 82 -811
rect 32 -814 103 -812
rect -68 -820 13 -815
rect -164 -863 -160 -859
rect -176 -867 -160 -863
rect -210 -888 -200 -883
rect -193 -884 -189 -871
rect -164 -879 -160 -867
rect -193 -889 -180 -884
rect -193 -891 -189 -889
rect -156 -864 -152 -859
rect -156 -868 -139 -864
rect -156 -879 -152 -868
rect -143 -878 -139 -868
rect -131 -878 -127 -866
rect -143 -883 -127 -878
rect -201 -950 -197 -911
rect -160 -931 -156 -918
rect -143 -944 -137 -883
rect -131 -886 -127 -883
rect -123 -879 -119 -866
rect -123 -883 -102 -879
rect -123 -886 -119 -883
rect -108 -884 -102 -883
rect -108 -889 -98 -884
rect -92 -889 -87 -884
rect -80 -885 -76 -872
rect -38 -846 -29 -833
rect 10 -840 13 -820
rect 45 -820 48 -814
rect 64 -820 67 -814
rect 79 -815 103 -814
rect 85 -821 88 -815
rect 54 -835 57 -832
rect 54 -838 67 -835
rect 10 -843 46 -840
rect 64 -841 67 -838
rect 64 -844 86 -841
rect 94 -841 97 -833
rect 94 -844 106 -841
rect -38 -849 56 -846
rect -80 -890 -63 -885
rect -80 -892 -76 -890
rect -127 -931 -123 -918
rect -88 -950 -84 -912
rect -38 -930 -30 -849
rect 64 -852 67 -844
rect 94 -847 97 -844
rect 995 -849 999 -810
rect 1036 -830 1040 -817
rect 1053 -840 1059 -782
rect 1065 -785 1069 -782
rect 1073 -778 1077 -765
rect 1387 -742 1400 -717
rect 1431 -742 1444 -717
rect 1316 -753 1333 -749
rect 1353 -750 1357 -742
rect 1353 -753 1393 -750
rect 1343 -761 1346 -757
rect 1353 -764 1357 -753
rect 1365 -761 1369 -756
rect 1389 -761 1393 -753
rect 1397 -756 1400 -742
rect 1441 -751 1444 -742
rect 1441 -756 1465 -751
rect 1472 -752 1476 -742
rect 1397 -761 1413 -756
rect 1433 -761 1437 -757
rect 1397 -764 1400 -761
rect 1441 -764 1444 -756
rect 1472 -757 1485 -752
rect 1472 -764 1476 -757
rect 1073 -782 1094 -778
rect 1073 -785 1077 -782
rect 1088 -783 1094 -782
rect 1088 -788 1098 -783
rect 1104 -788 1109 -783
rect 1116 -784 1120 -771
rect 1345 -774 1357 -764
rect 1389 -774 1400 -764
rect 1433 -774 1444 -764
rect 1333 -779 1337 -774
rect 1369 -779 1373 -774
rect 1413 -779 1417 -774
rect 1464 -779 1468 -774
rect 1332 -783 1476 -779
rect 1116 -789 1133 -784
rect 1116 -791 1120 -789
rect 1158 -792 1176 -786
rect 1069 -830 1073 -817
rect 1108 -849 1112 -811
rect 1158 -829 1166 -792
rect 85 -857 88 -853
rect 967 -857 1176 -849
rect 75 -860 103 -857
rect 45 -870 48 -864
rect 75 -870 79 -860
rect -20 -873 79 -870
rect -20 -950 -9 -873
rect -229 -951 -9 -950
rect -313 -958 -9 -951
<< m2contact >>
rect 985 166 991 171
rect -581 65 -570 72
rect -244 98 -238 103
rect -368 65 -357 72
rect -228 86 -223 91
rect -196 86 -191 91
rect -72 98 -62 105
rect 1001 154 1006 159
rect 1033 154 1038 159
rect 1085 154 1093 159
rect -144 86 -136 91
rect -283 18 -278 23
rect -248 17 -242 22
rect -228 -30 -223 -25
rect -107 73 -96 79
rect -166 17 -160 22
rect 946 86 951 91
rect 981 85 987 90
rect -131 16 -125 21
rect -195 -30 -190 -25
rect -106 -30 -98 -24
rect 285 44 291 49
rect 301 32 306 37
rect 333 32 338 37
rect 385 32 393 37
rect 246 -36 251 -31
rect 281 -37 287 -32
rect 215 -106 226 -97
rect 301 -84 306 -79
rect 493 26 498 32
rect 363 -37 369 -32
rect 398 -38 404 -33
rect 334 -84 339 -79
rect 318 -95 324 -90
rect 423 -84 431 -78
rect 493 -36 498 -30
rect 1001 38 1006 43
rect 1276 119 1281 124
rect 1063 85 1069 90
rect 1098 84 1104 89
rect 1034 38 1039 43
rect 1018 27 1024 33
rect 1123 38 1131 44
rect 482 -95 488 -90
rect 690 -91 695 -86
rect -566 -264 -555 -257
rect -229 -231 -223 -226
rect -353 -264 -342 -257
rect -213 -243 -208 -238
rect -181 -243 -176 -238
rect -57 -231 -47 -224
rect -129 -243 -121 -238
rect -268 -311 -263 -306
rect -233 -312 -227 -307
rect -213 -359 -208 -354
rect -92 -256 -81 -250
rect -151 -312 -145 -307
rect -116 -313 -110 -308
rect -180 -359 -175 -354
rect -91 -359 -83 -353
rect 280 -161 286 -156
rect 296 -173 301 -168
rect 328 -173 333 -168
rect 975 -142 981 -137
rect 380 -173 388 -168
rect 215 -251 220 -240
rect 241 -241 246 -236
rect 276 -242 282 -237
rect 296 -289 301 -284
rect 488 -179 493 -173
rect 358 -242 364 -237
rect 393 -243 399 -238
rect 329 -289 334 -284
rect 313 -300 319 -295
rect 418 -289 426 -283
rect 488 -241 493 -235
rect 991 -154 996 -149
rect 1023 -154 1028 -149
rect 1075 -154 1083 -149
rect 936 -222 941 -217
rect 971 -223 977 -218
rect 478 -270 483 -265
rect 477 -300 483 -295
rect 991 -270 996 -265
rect 1266 -189 1271 -184
rect 1053 -223 1059 -218
rect 1088 -224 1094 -219
rect 1024 -270 1029 -265
rect 1008 -281 1014 -275
rect 1113 -270 1121 -264
rect 688 -296 693 -291
rect 215 -317 222 -311
rect -542 -531 -531 -524
rect -205 -498 -199 -493
rect -329 -531 -318 -524
rect -189 -510 -184 -505
rect -157 -510 -152 -505
rect -33 -498 -23 -491
rect -105 -510 -97 -505
rect -244 -578 -239 -573
rect -209 -579 -203 -574
rect -189 -626 -184 -621
rect -68 -523 -57 -517
rect -127 -579 -121 -574
rect -92 -580 -86 -575
rect -156 -626 -151 -621
rect -67 -626 -59 -620
rect 329 -415 335 -410
rect 345 -427 350 -422
rect 377 -427 382 -422
rect 429 -427 437 -422
rect 290 -495 295 -490
rect 325 -496 331 -491
rect 255 -509 263 -498
rect 255 -565 270 -556
rect 345 -543 350 -538
rect 537 -433 542 -427
rect 407 -496 413 -491
rect 442 -497 448 -492
rect 378 -543 383 -538
rect 362 -554 368 -549
rect 467 -543 475 -537
rect 537 -495 542 -489
rect 518 -509 525 -500
rect 999 -401 1005 -396
rect 1015 -413 1020 -408
rect 1047 -413 1052 -408
rect 1099 -413 1107 -408
rect 960 -481 965 -476
rect 995 -482 1001 -477
rect 526 -554 532 -549
rect 1015 -529 1020 -524
rect 1290 -448 1295 -443
rect 1077 -482 1083 -477
rect 1112 -483 1118 -478
rect 1048 -529 1053 -524
rect 1032 -540 1038 -534
rect 1137 -529 1145 -523
rect 734 -550 739 -545
rect 324 -620 330 -615
rect 340 -632 345 -627
rect 372 -632 377 -627
rect 424 -632 432 -627
rect 259 -710 264 -699
rect 285 -700 290 -695
rect 320 -701 326 -696
rect 340 -748 345 -743
rect 532 -638 537 -632
rect 402 -701 408 -696
rect 437 -702 443 -697
rect 373 -748 378 -743
rect 357 -759 363 -754
rect 462 -748 470 -742
rect 532 -700 537 -694
rect 522 -729 527 -724
rect 521 -759 527 -754
rect 1020 -707 1026 -702
rect 1036 -719 1041 -714
rect 1068 -719 1073 -714
rect 1120 -719 1128 -714
rect 981 -787 986 -782
rect 1016 -788 1022 -783
rect -513 -841 -502 -834
rect -176 -808 -170 -803
rect -300 -841 -289 -834
rect -160 -820 -155 -815
rect -128 -820 -123 -815
rect -4 -808 6 -801
rect -76 -820 -68 -815
rect -215 -888 -210 -883
rect -180 -889 -174 -884
rect -160 -936 -155 -931
rect -39 -833 -28 -827
rect -98 -889 -92 -884
rect -63 -890 -57 -885
rect -127 -936 -122 -931
rect 1036 -835 1041 -830
rect 1311 -754 1316 -749
rect 1098 -788 1104 -783
rect 1133 -789 1139 -784
rect 1069 -835 1074 -830
rect 1053 -846 1059 -840
rect 1158 -835 1166 -829
rect -38 -936 -30 -930
<< metal2 >>
rect 991 166 1104 171
rect 946 154 1001 159
rect 1006 154 1033 159
rect 1038 154 1085 159
rect -342 134 -338 135
rect -342 130 -64 134
rect -555 119 -360 123
rect -555 71 -551 119
rect -570 66 -551 71
rect -342 71 -338 130
rect -299 121 -99 125
rect -238 98 -125 103
rect -357 66 -338 71
rect -283 86 -228 91
rect -223 86 -196 91
rect -191 86 -144 91
rect -283 23 -279 86
rect -248 -25 -242 17
rect -166 -24 -160 17
rect -131 21 -125 98
rect -105 79 -99 121
rect -69 105 -64 130
rect 946 91 950 154
rect 291 44 404 49
rect 246 32 301 37
rect 306 32 333 37
rect 338 32 385 37
rect -249 -30 -228 -25
rect -223 -30 -195 -25
rect -190 -30 -176 -25
rect -166 -30 -106 -24
rect 246 -31 250 32
rect 281 -79 287 -37
rect 363 -78 369 -37
rect 398 -33 404 44
rect 981 43 987 85
rect 1063 44 1069 85
rect 1098 89 1104 166
rect 980 38 1001 43
rect 1006 38 1034 43
rect 1039 38 1053 43
rect 1063 38 1123 44
rect 1276 31 1281 119
rect 1024 27 1281 31
rect 493 -30 498 26
rect 280 -84 301 -79
rect 306 -84 334 -79
rect 339 -84 353 -79
rect 363 -84 423 -78
rect 324 -95 482 -90
rect 690 -97 695 -91
rect 611 -103 695 -97
rect -327 -195 -323 -194
rect -327 -199 -49 -195
rect -540 -210 -345 -206
rect -540 -258 -536 -210
rect -555 -263 -536 -258
rect -327 -258 -323 -199
rect -284 -208 -84 -204
rect -223 -231 -110 -226
rect -342 -263 -323 -258
rect -268 -243 -213 -238
rect -208 -243 -181 -238
rect -176 -243 -129 -238
rect -268 -306 -264 -243
rect -233 -354 -227 -312
rect -151 -353 -145 -312
rect -116 -308 -110 -231
rect -90 -250 -84 -208
rect -54 -224 -49 -199
rect 215 -240 220 -106
rect 611 -126 617 -103
rect 473 -131 617 -126
rect 286 -161 399 -156
rect 241 -173 296 -168
rect 301 -173 328 -168
rect 333 -173 380 -168
rect 241 -236 245 -173
rect 276 -284 282 -242
rect 358 -283 364 -242
rect 393 -238 399 -161
rect 473 -270 478 -131
rect 981 -142 1094 -137
rect 936 -154 991 -149
rect 996 -154 1023 -149
rect 1028 -154 1075 -149
rect 488 -235 493 -179
rect 936 -217 940 -154
rect 971 -265 977 -223
rect 1053 -264 1059 -223
rect 1088 -219 1094 -142
rect 970 -270 991 -265
rect 996 -270 1024 -265
rect 1029 -270 1043 -265
rect 1053 -270 1113 -264
rect 1266 -277 1271 -189
rect 1014 -281 1271 -277
rect 275 -289 296 -284
rect 301 -289 329 -284
rect 334 -289 348 -284
rect 358 -289 418 -283
rect 319 -300 477 -295
rect -234 -359 -213 -354
rect -208 -359 -180 -354
rect -175 -359 -161 -354
rect -151 -359 -91 -353
rect -303 -462 -299 -461
rect -303 -466 -25 -462
rect -516 -477 -321 -473
rect -516 -525 -512 -477
rect -531 -530 -512 -525
rect -303 -525 -299 -466
rect -260 -475 -60 -471
rect -199 -498 -86 -493
rect -318 -530 -299 -525
rect -244 -510 -189 -505
rect -184 -510 -157 -505
rect -152 -510 -105 -505
rect -244 -573 -240 -510
rect -209 -621 -203 -579
rect -127 -620 -121 -579
rect -92 -575 -86 -498
rect -66 -517 -60 -475
rect -30 -491 -25 -466
rect 215 -491 222 -317
rect 688 -378 693 -296
rect 518 -384 693 -378
rect 335 -415 448 -410
rect 290 -427 345 -422
rect 350 -427 377 -422
rect 382 -427 429 -422
rect 290 -490 294 -427
rect 215 -498 263 -491
rect 325 -538 331 -496
rect 407 -537 413 -496
rect 442 -492 448 -415
rect 518 -500 525 -384
rect 1005 -401 1118 -396
rect 960 -413 1015 -408
rect 1020 -413 1047 -408
rect 1052 -413 1099 -408
rect 537 -489 542 -433
rect 960 -476 964 -413
rect 995 -524 1001 -482
rect 1077 -523 1083 -482
rect 1112 -478 1118 -401
rect 994 -529 1015 -524
rect 1020 -529 1048 -524
rect 1053 -529 1067 -524
rect 1077 -529 1137 -523
rect 324 -543 345 -538
rect 350 -543 378 -538
rect 383 -543 397 -538
rect 407 -543 467 -537
rect 1290 -536 1295 -448
rect 1038 -540 1295 -536
rect 368 -554 526 -549
rect 734 -556 739 -550
rect 655 -562 739 -556
rect -210 -626 -189 -621
rect -184 -626 -156 -621
rect -151 -626 -137 -621
rect -127 -626 -67 -620
rect 259 -699 264 -565
rect 655 -585 661 -562
rect 517 -590 661 -585
rect 330 -620 443 -615
rect 285 -632 340 -627
rect 345 -632 372 -627
rect 377 -632 424 -627
rect 285 -695 289 -632
rect 320 -743 326 -701
rect 402 -742 408 -701
rect 437 -697 443 -620
rect 517 -729 522 -590
rect 532 -694 537 -638
rect 1026 -707 1139 -702
rect 981 -719 1036 -714
rect 1041 -719 1068 -714
rect 1073 -719 1120 -714
rect 319 -748 340 -743
rect 345 -748 373 -743
rect 378 -748 392 -743
rect 402 -748 462 -742
rect 363 -759 521 -754
rect -274 -772 -270 -771
rect -274 -776 4 -772
rect -487 -787 -292 -783
rect -487 -835 -483 -787
rect -502 -840 -483 -835
rect -274 -835 -270 -776
rect -231 -785 -31 -781
rect -170 -808 -57 -803
rect -289 -840 -270 -835
rect -215 -820 -160 -815
rect -155 -820 -128 -815
rect -123 -820 -76 -815
rect -215 -883 -211 -820
rect -180 -931 -174 -889
rect -98 -930 -92 -889
rect -63 -885 -57 -808
rect -37 -827 -31 -785
rect -1 -801 4 -776
rect 981 -782 985 -719
rect 1016 -830 1022 -788
rect 1098 -829 1104 -788
rect 1133 -784 1139 -707
rect 1015 -835 1036 -830
rect 1041 -835 1069 -830
rect 1074 -835 1088 -830
rect 1098 -835 1158 -829
rect 1311 -842 1316 -754
rect 1059 -846 1316 -842
rect -181 -936 -160 -931
rect -155 -936 -127 -931
rect -122 -936 -108 -931
rect -98 -936 -38 -930
<< m3contact >>
rect -360 118 -347 124
rect -309 119 -299 125
rect -345 -211 -332 -205
rect -294 -210 -284 -204
rect -321 -478 -308 -472
rect -270 -477 -260 -471
rect -292 -788 -279 -782
rect -241 -787 -231 -781
<< metal3 >>
rect -347 119 -309 124
rect -332 -210 -294 -205
rect -308 -477 -270 -472
rect -279 -787 -241 -782
<< labels >>
rlabel metal1 457 32 472 37 1 a0_reg
rlabel metal1 423 -19 431 -3 1 b0_reg
rlabel metal1 341 57 455 62 1 vdd
rlabel metal1 317 -105 431 -99 1 gnd
rlabel metal1 318 -90 324 -85 1 p0
rlabel metal1 336 -148 450 -143 1 vdd
rlabel metal1 675 -260 675 -260 1 gnd!
rlabel metal1 312 -310 426 -304 1 gnd
rlabel metal1 313 -295 319 -290 1 p1
rlabel metal1 418 -224 426 -208 1 b1_reg
rlabel metal1 452 -173 467 -168 1 a1_reg
rlabel metal1 673 -245 679 -242 1 c1
rlabel metal1 678 -40 684 -37 1 c0
rlabel metal1 356 -769 470 -763 1 gnd
rlabel metal1 676 -661 676 -661 5 vdd!
rlabel metal1 679 -726 679 -726 1 gnd!
rlabel metal1 713 -674 713 -674 5 vdd!
rlabel metal1 719 -719 719 -719 1 gnd!
rlabel metal1 380 -607 494 -602 1 vdd
rlabel metal1 724 -514 724 -514 1 gnd!
rlabel metal1 718 -469 718 -469 5 vdd!
rlabel metal1 684 -521 684 -521 1 gnd!
rlabel metal1 681 -456 681 -456 5 vdd!
rlabel metal1 361 -564 475 -558 1 gnd
rlabel metal1 385 -402 499 -397 1 vdd
rlabel metal1 362 -549 368 -544 1 p2
rlabel metal1 467 -478 475 -462 1 b2_reg
rlabel metal1 501 -427 516 -422 1 a2_reg
rlabel metal1 357 -754 363 -749 1 p3
rlabel metal1 496 -632 511 -627 1 a3_reg
rlabel metal1 462 -683 470 -667 1 b3_reg
rlabel metal1 717 -704 723 -701 1 out_carry
rlabel metal1 722 -499 728 -496 1 c2
rlabel metal1 -211 -37 -205 -31 1 p0
rlabel metal1 -188 111 -74 116 1 vdd
rlabel metal1 -212 -51 -98 -45 1 gnd
rlabel metal1 -510 63 -508 65 1 clk
rlabel metal1 -512 42 -509 43 1 gnd
rlabel metal1 -506 114 -504 115 5 vdd
rlabel metal1 -487 63 -486 65 1 clk
rlabel metal1 -419 63 -417 65 1 clk
rlabel metal1 -375 68 -372 70 1 a0_reg
rlabel metal1 -525 71 -523 73 3 a0
rlabel metal1 -632 63 -630 65 1 clk
rlabel metal1 -700 63 -699 65 1 clk
rlabel metal1 -719 114 -717 115 5 vdd
rlabel metal1 -725 42 -722 43 1 gnd
rlabel metal1 -723 63 -721 65 1 clk
rlabel metal1 -738 71 -736 73 3 b0
rlabel metal1 -588 68 -585 70 1 b0_reg
rlabel metal1 -173 -218 -59 -213 1 vdd
rlabel metal1 -197 -380 -83 -374 1 gnd
rlabel metal1 -495 -266 -493 -264 1 clk
rlabel metal1 -497 -287 -494 -286 1 gnd
rlabel metal1 -491 -215 -489 -214 5 vdd
rlabel metal1 -472 -266 -471 -264 1 clk
rlabel metal1 -404 -266 -402 -264 1 clk
rlabel metal1 -617 -266 -615 -264 1 clk
rlabel metal1 -685 -266 -684 -264 1 clk
rlabel metal1 -704 -215 -702 -214 5 vdd
rlabel metal1 -710 -287 -707 -286 1 gnd
rlabel metal1 -708 -266 -706 -264 1 clk
rlabel metal1 70 -549 70 -549 1 gnd!
rlabel metal1 -149 -485 -35 -480 1 vdd
rlabel metal1 -173 -647 -59 -641 1 gnd
rlabel metal1 -471 -533 -469 -531 1 clk
rlabel metal1 -473 -554 -470 -553 1 gnd
rlabel metal1 -467 -482 -465 -481 5 vdd
rlabel metal1 -448 -533 -447 -531 1 clk
rlabel metal1 -380 -533 -378 -531 1 clk
rlabel metal1 -593 -533 -591 -531 1 clk
rlabel metal1 -661 -533 -660 -531 1 clk
rlabel metal1 -680 -482 -678 -481 5 vdd
rlabel metal1 -686 -554 -683 -553 1 gnd
rlabel metal1 -684 -533 -682 -531 1 clk
rlabel metal1 -655 -843 -653 -841 1 clk
rlabel metal1 -657 -864 -654 -863 1 gnd
rlabel metal1 -651 -792 -649 -791 5 vdd
rlabel metal1 -632 -843 -631 -841 1 clk
rlabel metal1 -564 -843 -562 -841 1 clk
rlabel metal1 -351 -843 -349 -841 1 clk
rlabel metal1 -419 -843 -418 -841 1 clk
rlabel metal1 -438 -792 -436 -791 5 vdd
rlabel metal1 -444 -864 -441 -863 1 gnd
rlabel metal1 -442 -843 -440 -841 1 clk
rlabel metal1 -144 -957 -30 -951 1 gnd
rlabel metal1 -120 -795 -6 -790 1 vdd
rlabel metal1 99 -859 99 -859 1 gnd!
rlabel metal1 -510 -258 -508 -256 1 a1
rlabel metal1 -575 -261 -570 -259 1 b1_reg
rlabel metal1 -723 -258 -721 -256 1 b1
rlabel metal1 -360 -261 -357 -259 1 a1_reg
rlabel metal1 -196 -366 -190 -360 1 p1
rlabel metal1 -57 -243 -42 -238 1 a1_reg
rlabel metal1 48 -267 53 -264 1 g1
rlabel metal1 -486 -525 -484 -523 1 a2
rlabel metal1 -336 -528 -333 -526 1 a2_reg
rlabel metal1 -549 -528 -546 -526 1 b2_reg
rlabel metal1 -699 -525 -696 -523 1 b2
rlabel metal1 -172 -633 -166 -627 1 p2
rlabel metal1 72 -534 77 -531 1 g2
rlabel metal1 101 -844 106 -841 7 g3
rlabel metal1 -91 -294 -83 -277 1 b1_reg
rlabel metal1 -143 -943 -137 -937 1 p3
rlabel metal1 -307 -838 -304 -836 1 a3_reg
rlabel metal1 -457 -835 -454 -833 1 a3
rlabel metal1 -520 -838 -517 -836 1 b3_reg
rlabel metal1 -670 -835 -667 -833 1 b3
rlabel metal1 1017 17 1131 23 1 GND
rlabel metal1 1041 179 1155 184 5 VDD
rlabel metal1 1123 81 1139 87 1 p0
rlabel metal1 1399 113 1401 115 1 clk
rlabel metal1 1331 113 1332 115 1 clk
rlabel metal1 1312 164 1314 165 5 vdd
rlabel metal1 1306 92 1309 93 1 gnd
rlabel metal1 1308 113 1310 115 1 clk
rlabel metal1 1443 118 1446 120 1 s0_reg
rlabel metal1 1293 121 1295 123 1 s0
rlabel metal1 1018 34 1024 38 1 s0
rlabel metal1 1007 -291 1121 -285 1 GND
rlabel metal1 1031 -129 1145 -124 5 VDD
rlabel metal1 1389 -195 1391 -193 1 clk
rlabel metal1 1321 -195 1322 -193 1 clk
rlabel metal1 1302 -144 1304 -143 5 vdd
rlabel metal1 1296 -216 1299 -215 1 gnd
rlabel metal1 1298 -195 1300 -193 1 clk
rlabel metal1 1031 -550 1145 -544 1 GND
rlabel metal1 1055 -388 1169 -383 5 VDD
rlabel metal1 1413 -454 1415 -452 1 clk
rlabel metal1 1345 -454 1346 -452 1 clk
rlabel metal1 1326 -403 1328 -402 5 vdd
rlabel metal1 1320 -475 1323 -474 1 gnd
rlabel metal1 1322 -454 1324 -452 1 clk
rlabel metal1 1052 -856 1166 -850 1 GND
rlabel metal1 1076 -694 1190 -689 5 VDD
rlabel metal1 1434 -760 1436 -758 1 clk
rlabel metal1 1366 -760 1367 -758 1 clk
rlabel metal1 1347 -709 1349 -708 5 vdd
rlabel metal1 1341 -781 1344 -780 1 gnd
rlabel metal1 1343 -760 1345 -758 1 clk
rlabel metal1 1283 -187 1285 -185 1 s1
rlabel metal1 1433 -190 1436 -188 1 s1_reg
rlabel metal1 1008 -274 1014 -270 1 s1
rlabel metal1 1032 -533 1038 -529 1 s2
rlabel metal1 1053 -839 1059 -835 1 s3
rlabel metal1 1307 -446 1309 -444 1 s2
rlabel metal1 1457 -449 1460 -447 1 s2_reg
rlabel metal1 1478 -755 1481 -753 1 s3_reg
rlabel metal1 1328 -752 1330 -750 1 s3
rlabel metal1 1119 -148 1156 -143 1 c0
rlabel metal1 1113 -227 1129 -221 1 p1
rlabel metal1 1137 -486 1153 -480 1 p2
rlabel metal1 1143 -407 1180 -402 1 c1
rlabel metal1 1158 -792 1174 -786 1 p3
rlabel metal1 1164 -713 1201 -708 1 c2
rlabel metal1 1129 160 1166 165 1 carry_reg
rlabel metal1 698 58 700 60 1 clk
rlabel metal1 696 37 699 38 1 gnd
rlabel metal1 702 109 704 110 5 vdd
rlabel metal1 721 58 722 60 1 clk
rlabel metal1 789 58 791 60 1 clk
rlabel metal1 832 63 837 65 1 carry_reg
rlabel metal1 683 66 685 68 3 carry
rlabel metal1 33 62 38 65 1 g0
rlabel metal1 505 -65 509 -62 1 carry_reg
rlabel metal1 632 -202 632 -202 5 vdd!
rlabel metal1 635 -267 635 -267 1 gnd!
rlabel metal1 669 -215 669 -215 5 vdd!
rlabel metal1 505 -71 508 -68 1 p0
rlabel metal1 885 -715 890 -713 1 out_carry_reg
rlabel metal1 842 -720 844 -718 1 clk
rlabel metal1 774 -720 775 -718 1 clk
rlabel metal1 755 -669 757 -668 5 vdd
rlabel metal1 749 -741 752 -740 1 gnd
rlabel metal1 751 -720 753 -718 1 clk
<< end >>
