magic
tech scmos
timestamp 1618579805
<< nwell >>
rect 0 6 24 30
<< polysilicon >>
rect 11 24 13 27
rect 11 -2 13 12
rect 11 -11 13 -8
<< ndiffusion >>
rect 10 -8 11 -2
rect 13 -8 14 -2
<< pdiffusion >>
rect 10 12 11 24
rect 13 12 14 24
<< metal1 >>
rect 0 30 24 33
rect 6 24 9 30
rect 0 1 7 4
rect 15 4 18 12
rect 15 1 24 4
rect 15 -2 18 1
rect 6 -12 9 -8
rect 0 -15 24 -12
<< ntransistor >>
rect 11 -8 13 -2
<< ptransistor >>
rect 11 12 13 24
<< polycontact >>
rect 7 1 11 5
<< ndcontact >>
rect 6 -8 10 -2
rect 14 -8 18 -2
<< pdcontact >>
rect 6 12 10 24
rect 14 12 18 24
<< labels >>
rlabel metal1 14 31 14 31 5 vdd!
rlabel metal1 20 -14 20 -14 1 gnd!
rlabel metal1 0 1 0 4 3 in
rlabel metal1 24 1 24 4 7 op
<< end >>
