magic
tech scmos
timestamp 1731738108
<< nwell >>
rect -205 39 -173 76
rect -167 39 -141 76
rect -123 39 -97 76
rect -78 39 -52 76
rect 8 39 40 76
rect 46 39 72 76
rect 90 39 116 76
rect 135 39 161 76
rect 255 -11 280 46
rect 292 -39 317 1
rect 325 -6 350 34
rect 368 -12 393 45
rect 501 32 535 56
rect 541 31 565 55
rect -190 -290 -158 -253
rect -152 -290 -126 -253
rect -108 -290 -82 -253
rect -63 -290 -37 -253
rect 23 -290 55 -253
rect 61 -290 87 -253
rect 105 -290 131 -253
rect 150 -290 176 -253
rect 270 -340 295 -283
rect 307 -368 332 -328
rect 340 -335 365 -295
rect 383 -341 408 -284
rect 516 -297 550 -273
rect 556 -298 580 -274
rect -166 -557 -134 -520
rect -128 -557 -102 -520
rect -84 -557 -58 -520
rect -39 -557 -13 -520
rect 47 -557 79 -520
rect 85 -557 111 -520
rect 129 -557 155 -520
rect 174 -557 200 -520
rect 294 -607 319 -550
rect 331 -635 356 -595
rect 364 -602 389 -562
rect 407 -608 432 -551
rect 540 -564 574 -540
rect 580 -565 604 -541
rect -137 -867 -105 -830
rect -99 -867 -73 -830
rect -55 -867 -29 -830
rect -10 -867 16 -830
rect 76 -867 108 -830
rect 114 -867 140 -830
rect 158 -867 184 -830
rect 203 -867 229 -830
rect 323 -917 348 -860
rect 360 -945 385 -905
rect 393 -912 418 -872
rect 436 -918 461 -861
rect 569 -874 603 -850
rect 609 -875 633 -851
<< ntransistor >>
rect -198 13 -196 23
rect -162 13 -160 23
rect -154 13 -152 23
rect -118 13 -116 23
rect -110 13 -108 23
rect -67 13 -65 23
rect 15 13 17 23
rect 51 13 53 23
rect 59 13 61 23
rect 95 13 97 23
rect 103 13 105 23
rect 146 13 148 23
rect 303 11 305 31
rect 512 6 514 18
rect 522 6 524 18
rect 552 17 554 23
rect 266 -41 268 -21
rect 336 -36 338 -16
rect 379 -42 381 -22
rect -183 -316 -181 -306
rect -147 -316 -145 -306
rect -139 -316 -137 -306
rect -103 -316 -101 -306
rect -95 -316 -93 -306
rect -52 -316 -50 -306
rect 30 -316 32 -306
rect 66 -316 68 -306
rect 74 -316 76 -306
rect 110 -316 112 -306
rect 118 -316 120 -306
rect 161 -316 163 -306
rect 318 -318 320 -298
rect 527 -323 529 -311
rect 537 -323 539 -311
rect 567 -312 569 -306
rect 281 -370 283 -350
rect 351 -365 353 -345
rect 394 -371 396 -351
rect -159 -583 -157 -573
rect -123 -583 -121 -573
rect -115 -583 -113 -573
rect -79 -583 -77 -573
rect -71 -583 -69 -573
rect -28 -583 -26 -573
rect 54 -583 56 -573
rect 90 -583 92 -573
rect 98 -583 100 -573
rect 134 -583 136 -573
rect 142 -583 144 -573
rect 185 -583 187 -573
rect 342 -585 344 -565
rect 551 -590 553 -578
rect 561 -590 563 -578
rect 591 -579 593 -573
rect 305 -637 307 -617
rect 375 -632 377 -612
rect 418 -638 420 -618
rect -130 -893 -128 -883
rect -94 -893 -92 -883
rect -86 -893 -84 -883
rect -50 -893 -48 -883
rect -42 -893 -40 -883
rect 1 -893 3 -883
rect 83 -893 85 -883
rect 119 -893 121 -883
rect 127 -893 129 -883
rect 163 -893 165 -883
rect 171 -893 173 -883
rect 214 -893 216 -883
rect 371 -895 373 -875
rect 580 -900 582 -888
rect 590 -900 592 -888
rect 620 -889 622 -883
rect 334 -947 336 -927
rect 404 -942 406 -922
rect 447 -948 449 -928
<< ptransistor >>
rect -194 45 -192 70
rect -186 45 -184 70
rect -156 45 -154 70
rect -112 45 -110 70
rect -67 45 -65 70
rect 19 45 21 70
rect 27 45 29 70
rect 57 45 59 70
rect 101 45 103 70
rect 146 45 148 70
rect 266 -1 268 39
rect 512 38 514 50
rect 522 38 524 50
rect 336 4 338 24
rect 379 -2 381 38
rect 552 37 554 49
rect 303 -29 305 -9
rect -179 -284 -177 -259
rect -171 -284 -169 -259
rect -141 -284 -139 -259
rect -97 -284 -95 -259
rect -52 -284 -50 -259
rect 34 -284 36 -259
rect 42 -284 44 -259
rect 72 -284 74 -259
rect 116 -284 118 -259
rect 161 -284 163 -259
rect 281 -330 283 -290
rect 527 -291 529 -279
rect 537 -291 539 -279
rect 351 -325 353 -305
rect 394 -331 396 -291
rect 567 -292 569 -280
rect 318 -358 320 -338
rect -155 -551 -153 -526
rect -147 -551 -145 -526
rect -117 -551 -115 -526
rect -73 -551 -71 -526
rect -28 -551 -26 -526
rect 58 -551 60 -526
rect 66 -551 68 -526
rect 96 -551 98 -526
rect 140 -551 142 -526
rect 185 -551 187 -526
rect 305 -597 307 -557
rect 551 -558 553 -546
rect 561 -558 563 -546
rect 375 -592 377 -572
rect 418 -598 420 -558
rect 591 -559 593 -547
rect 342 -625 344 -605
rect -126 -861 -124 -836
rect -118 -861 -116 -836
rect -88 -861 -86 -836
rect -44 -861 -42 -836
rect 1 -861 3 -836
rect 87 -861 89 -836
rect 95 -861 97 -836
rect 125 -861 127 -836
rect 169 -861 171 -836
rect 214 -861 216 -836
rect 334 -907 336 -867
rect 580 -868 582 -856
rect 590 -868 592 -856
rect 404 -902 406 -882
rect 447 -908 449 -868
rect 620 -869 622 -857
rect 371 -935 373 -915
<< ndiffusion >>
rect -199 13 -198 23
rect -196 13 -195 23
rect -163 13 -162 23
rect -160 13 -159 23
rect -155 13 -154 23
rect -152 13 -151 23
rect -119 13 -118 23
rect -116 13 -115 23
rect -111 13 -110 23
rect -108 13 -107 23
rect -68 13 -67 23
rect -65 13 -64 23
rect 14 13 15 23
rect 17 13 18 23
rect 50 13 51 23
rect 53 13 54 23
rect 58 13 59 23
rect 61 13 62 23
rect 94 13 95 23
rect 97 13 98 23
rect 102 13 103 23
rect 105 13 106 23
rect 145 13 146 23
rect 148 13 149 23
rect 302 11 303 31
rect 305 11 306 31
rect 511 6 512 18
rect 514 6 522 18
rect 524 6 525 18
rect 551 17 552 23
rect 554 17 555 23
rect 265 -41 266 -21
rect 268 -41 269 -21
rect 335 -36 336 -16
rect 338 -36 339 -16
rect 378 -42 379 -22
rect 381 -42 382 -22
rect -184 -316 -183 -306
rect -181 -316 -180 -306
rect -148 -316 -147 -306
rect -145 -316 -144 -306
rect -140 -316 -139 -306
rect -137 -316 -136 -306
rect -104 -316 -103 -306
rect -101 -316 -100 -306
rect -96 -316 -95 -306
rect -93 -316 -92 -306
rect -53 -316 -52 -306
rect -50 -316 -49 -306
rect 29 -316 30 -306
rect 32 -316 33 -306
rect 65 -316 66 -306
rect 68 -316 69 -306
rect 73 -316 74 -306
rect 76 -316 77 -306
rect 109 -316 110 -306
rect 112 -316 113 -306
rect 117 -316 118 -306
rect 120 -316 121 -306
rect 160 -316 161 -306
rect 163 -316 164 -306
rect 317 -318 318 -298
rect 320 -318 321 -298
rect 526 -323 527 -311
rect 529 -323 537 -311
rect 539 -323 540 -311
rect 566 -312 567 -306
rect 569 -312 570 -306
rect 280 -370 281 -350
rect 283 -370 284 -350
rect 350 -365 351 -345
rect 353 -365 354 -345
rect 393 -371 394 -351
rect 396 -371 397 -351
rect -160 -583 -159 -573
rect -157 -583 -156 -573
rect -124 -583 -123 -573
rect -121 -583 -120 -573
rect -116 -583 -115 -573
rect -113 -583 -112 -573
rect -80 -583 -79 -573
rect -77 -583 -76 -573
rect -72 -583 -71 -573
rect -69 -583 -68 -573
rect -29 -583 -28 -573
rect -26 -583 -25 -573
rect 53 -583 54 -573
rect 56 -583 57 -573
rect 89 -583 90 -573
rect 92 -583 93 -573
rect 97 -583 98 -573
rect 100 -583 101 -573
rect 133 -583 134 -573
rect 136 -583 137 -573
rect 141 -583 142 -573
rect 144 -583 145 -573
rect 184 -583 185 -573
rect 187 -583 188 -573
rect 341 -585 342 -565
rect 344 -585 345 -565
rect 550 -590 551 -578
rect 553 -590 561 -578
rect 563 -590 564 -578
rect 590 -579 591 -573
rect 593 -579 594 -573
rect 304 -637 305 -617
rect 307 -637 308 -617
rect 374 -632 375 -612
rect 377 -632 378 -612
rect 417 -638 418 -618
rect 420 -638 421 -618
rect -131 -893 -130 -883
rect -128 -893 -127 -883
rect -95 -893 -94 -883
rect -92 -893 -91 -883
rect -87 -893 -86 -883
rect -84 -893 -83 -883
rect -51 -893 -50 -883
rect -48 -893 -47 -883
rect -43 -893 -42 -883
rect -40 -893 -39 -883
rect 0 -893 1 -883
rect 3 -893 4 -883
rect 82 -893 83 -883
rect 85 -893 86 -883
rect 118 -893 119 -883
rect 121 -893 122 -883
rect 126 -893 127 -883
rect 129 -893 130 -883
rect 162 -893 163 -883
rect 165 -893 166 -883
rect 170 -893 171 -883
rect 173 -893 174 -883
rect 213 -893 214 -883
rect 216 -893 217 -883
rect 370 -895 371 -875
rect 373 -895 374 -875
rect 579 -900 580 -888
rect 582 -900 590 -888
rect 592 -900 593 -888
rect 619 -889 620 -883
rect 622 -889 623 -883
rect 333 -947 334 -927
rect 336 -947 337 -927
rect 403 -942 404 -922
rect 406 -942 407 -922
rect 446 -948 447 -928
rect 449 -948 450 -928
<< pdiffusion >>
rect -195 45 -194 70
rect -192 45 -191 70
rect -187 45 -186 70
rect -184 45 -183 70
rect -157 45 -156 70
rect -154 45 -153 70
rect -113 45 -112 70
rect -110 45 -109 70
rect -68 45 -67 70
rect -65 45 -64 70
rect 18 45 19 70
rect 21 45 22 70
rect 26 45 27 70
rect 29 45 30 70
rect 56 45 57 70
rect 59 45 60 70
rect 100 45 101 70
rect 103 45 104 70
rect 145 45 146 70
rect 148 45 149 70
rect 265 -1 266 39
rect 268 -1 269 39
rect 511 38 512 50
rect 514 38 516 50
rect 520 38 522 50
rect 524 38 525 50
rect 335 4 336 24
rect 338 4 339 24
rect 378 -2 379 38
rect 381 -2 382 38
rect 551 37 552 49
rect 554 37 555 49
rect 302 -29 303 -9
rect 305 -29 306 -9
rect -180 -284 -179 -259
rect -177 -284 -176 -259
rect -172 -284 -171 -259
rect -169 -284 -168 -259
rect -142 -284 -141 -259
rect -139 -284 -138 -259
rect -98 -284 -97 -259
rect -95 -284 -94 -259
rect -53 -284 -52 -259
rect -50 -284 -49 -259
rect 33 -284 34 -259
rect 36 -284 37 -259
rect 41 -284 42 -259
rect 44 -284 45 -259
rect 71 -284 72 -259
rect 74 -284 75 -259
rect 115 -284 116 -259
rect 118 -284 119 -259
rect 160 -284 161 -259
rect 163 -284 164 -259
rect 280 -330 281 -290
rect 283 -330 284 -290
rect 526 -291 527 -279
rect 529 -291 531 -279
rect 535 -291 537 -279
rect 539 -291 540 -279
rect 350 -325 351 -305
rect 353 -325 354 -305
rect 393 -331 394 -291
rect 396 -331 397 -291
rect 566 -292 567 -280
rect 569 -292 570 -280
rect 317 -358 318 -338
rect 320 -358 321 -338
rect -156 -551 -155 -526
rect -153 -551 -152 -526
rect -148 -551 -147 -526
rect -145 -551 -144 -526
rect -118 -551 -117 -526
rect -115 -551 -114 -526
rect -74 -551 -73 -526
rect -71 -551 -70 -526
rect -29 -551 -28 -526
rect -26 -551 -25 -526
rect 57 -551 58 -526
rect 60 -551 61 -526
rect 65 -551 66 -526
rect 68 -551 69 -526
rect 95 -551 96 -526
rect 98 -551 99 -526
rect 139 -551 140 -526
rect 142 -551 143 -526
rect 184 -551 185 -526
rect 187 -551 188 -526
rect 304 -597 305 -557
rect 307 -597 308 -557
rect 550 -558 551 -546
rect 553 -558 555 -546
rect 559 -558 561 -546
rect 563 -558 564 -546
rect 374 -592 375 -572
rect 377 -592 378 -572
rect 417 -598 418 -558
rect 420 -598 421 -558
rect 590 -559 591 -547
rect 593 -559 594 -547
rect 341 -625 342 -605
rect 344 -625 345 -605
rect -127 -861 -126 -836
rect -124 -861 -123 -836
rect -119 -861 -118 -836
rect -116 -861 -115 -836
rect -89 -861 -88 -836
rect -86 -861 -85 -836
rect -45 -861 -44 -836
rect -42 -861 -41 -836
rect 0 -861 1 -836
rect 3 -861 4 -836
rect 86 -861 87 -836
rect 89 -861 90 -836
rect 94 -861 95 -836
rect 97 -861 98 -836
rect 124 -861 125 -836
rect 127 -861 128 -836
rect 168 -861 169 -836
rect 171 -861 172 -836
rect 213 -861 214 -836
rect 216 -861 217 -836
rect 333 -907 334 -867
rect 336 -907 337 -867
rect 579 -868 580 -856
rect 582 -868 584 -856
rect 588 -868 590 -856
rect 592 -868 593 -856
rect 403 -902 404 -882
rect 406 -902 407 -882
rect 446 -908 447 -868
rect 449 -908 450 -868
rect 619 -869 620 -857
rect 622 -869 623 -857
rect 370 -935 371 -915
rect 373 -935 374 -915
<< ndcontact >>
rect -203 13 -199 23
rect -195 13 -191 23
rect -167 13 -163 23
rect -159 13 -155 23
rect -151 13 -147 23
rect -123 13 -119 23
rect -115 13 -111 23
rect -107 13 -103 23
rect -72 13 -68 23
rect -64 13 -60 23
rect 10 13 14 23
rect 18 13 22 23
rect 46 13 50 23
rect 54 13 58 23
rect 62 13 66 23
rect 90 13 94 23
rect 98 13 102 23
rect 106 13 110 23
rect 141 13 145 23
rect 149 13 153 23
rect 298 11 302 31
rect 306 11 310 31
rect 507 6 511 18
rect 525 6 529 18
rect 547 17 551 23
rect 555 17 559 23
rect 261 -41 265 -21
rect 269 -41 273 -21
rect 331 -36 335 -16
rect 339 -36 343 -16
rect 374 -42 378 -22
rect 382 -42 386 -22
rect -188 -316 -184 -306
rect -180 -316 -176 -306
rect -152 -316 -148 -306
rect -144 -316 -140 -306
rect -136 -316 -132 -306
rect -108 -316 -104 -306
rect -100 -316 -96 -306
rect -92 -316 -88 -306
rect -57 -316 -53 -306
rect -49 -316 -45 -306
rect 25 -316 29 -306
rect 33 -316 37 -306
rect 61 -316 65 -306
rect 69 -316 73 -306
rect 77 -316 81 -306
rect 105 -316 109 -306
rect 113 -316 117 -306
rect 121 -316 125 -306
rect 156 -316 160 -306
rect 164 -316 168 -306
rect 313 -318 317 -298
rect 321 -318 325 -298
rect 522 -323 526 -311
rect 540 -323 544 -311
rect 562 -312 566 -306
rect 570 -312 574 -306
rect 276 -370 280 -350
rect 284 -370 288 -350
rect 346 -365 350 -345
rect 354 -365 358 -345
rect 389 -371 393 -351
rect 397 -371 401 -351
rect -164 -583 -160 -573
rect -156 -583 -152 -573
rect -128 -583 -124 -573
rect -120 -583 -116 -573
rect -112 -583 -108 -573
rect -84 -583 -80 -573
rect -76 -583 -72 -573
rect -68 -583 -64 -573
rect -33 -583 -29 -573
rect -25 -583 -21 -573
rect 49 -583 53 -573
rect 57 -583 61 -573
rect 85 -583 89 -573
rect 93 -583 97 -573
rect 101 -583 105 -573
rect 129 -583 133 -573
rect 137 -583 141 -573
rect 145 -583 149 -573
rect 180 -583 184 -573
rect 188 -583 192 -573
rect 337 -585 341 -565
rect 345 -585 349 -565
rect 546 -590 550 -578
rect 564 -590 568 -578
rect 586 -579 590 -573
rect 594 -579 598 -573
rect 300 -637 304 -617
rect 308 -637 312 -617
rect 370 -632 374 -612
rect 378 -632 382 -612
rect 413 -638 417 -618
rect 421 -638 425 -618
rect -135 -893 -131 -883
rect -127 -893 -123 -883
rect -99 -893 -95 -883
rect -91 -893 -87 -883
rect -83 -893 -79 -883
rect -55 -893 -51 -883
rect -47 -893 -43 -883
rect -39 -893 -35 -883
rect -4 -893 0 -883
rect 4 -893 8 -883
rect 78 -893 82 -883
rect 86 -893 90 -883
rect 114 -893 118 -883
rect 122 -893 126 -883
rect 130 -893 134 -883
rect 158 -893 162 -883
rect 166 -893 170 -883
rect 174 -893 178 -883
rect 209 -893 213 -883
rect 217 -893 221 -883
rect 366 -895 370 -875
rect 374 -895 378 -875
rect 575 -900 579 -888
rect 593 -900 597 -888
rect 615 -889 619 -883
rect 623 -889 627 -883
rect 329 -947 333 -927
rect 337 -947 341 -927
rect 399 -942 403 -922
rect 407 -942 411 -922
rect 442 -948 446 -928
rect 450 -948 454 -928
<< pdcontact >>
rect -199 45 -195 70
rect -191 45 -187 70
rect -183 45 -179 70
rect -161 45 -157 70
rect -153 45 -149 70
rect -117 45 -113 70
rect -109 45 -105 70
rect -72 45 -68 70
rect -64 45 -60 70
rect 14 45 18 70
rect 22 45 26 70
rect 30 45 34 70
rect 52 45 56 70
rect 60 45 64 70
rect 96 45 100 70
rect 104 45 108 70
rect 141 45 145 70
rect 149 45 153 70
rect 261 -1 265 39
rect 269 -1 273 39
rect 507 38 511 50
rect 516 38 520 50
rect 525 38 529 50
rect 331 4 335 24
rect 339 4 343 24
rect 374 -2 378 38
rect 382 -2 386 38
rect 547 37 551 49
rect 555 37 559 49
rect 298 -29 302 -9
rect 306 -29 310 -9
rect -184 -284 -180 -259
rect -176 -284 -172 -259
rect -168 -284 -164 -259
rect -146 -284 -142 -259
rect -138 -284 -134 -259
rect -102 -284 -98 -259
rect -94 -284 -90 -259
rect -57 -284 -53 -259
rect -49 -284 -45 -259
rect 29 -284 33 -259
rect 37 -284 41 -259
rect 45 -284 49 -259
rect 67 -284 71 -259
rect 75 -284 79 -259
rect 111 -284 115 -259
rect 119 -284 123 -259
rect 156 -284 160 -259
rect 164 -284 168 -259
rect 276 -330 280 -290
rect 284 -330 288 -290
rect 522 -291 526 -279
rect 531 -291 535 -279
rect 540 -291 544 -279
rect 346 -325 350 -305
rect 354 -325 358 -305
rect 389 -331 393 -291
rect 397 -331 401 -291
rect 562 -292 566 -280
rect 570 -292 574 -280
rect 313 -358 317 -338
rect 321 -358 325 -338
rect -160 -551 -156 -526
rect -152 -551 -148 -526
rect -144 -551 -140 -526
rect -122 -551 -118 -526
rect -114 -551 -110 -526
rect -78 -551 -74 -526
rect -70 -551 -66 -526
rect -33 -551 -29 -526
rect -25 -551 -21 -526
rect 53 -551 57 -526
rect 61 -551 65 -526
rect 69 -551 73 -526
rect 91 -551 95 -526
rect 99 -551 103 -526
rect 135 -551 139 -526
rect 143 -551 147 -526
rect 180 -551 184 -526
rect 188 -551 192 -526
rect 300 -597 304 -557
rect 308 -597 312 -557
rect 546 -558 550 -546
rect 555 -558 559 -546
rect 564 -558 568 -546
rect 370 -592 374 -572
rect 378 -592 382 -572
rect 413 -598 417 -558
rect 421 -598 425 -558
rect 586 -559 590 -547
rect 594 -559 598 -547
rect 337 -625 341 -605
rect 345 -625 349 -605
rect -131 -861 -127 -836
rect -123 -861 -119 -836
rect -115 -861 -111 -836
rect -93 -861 -89 -836
rect -85 -861 -81 -836
rect -49 -861 -45 -836
rect -41 -861 -37 -836
rect -4 -861 0 -836
rect 4 -861 8 -836
rect 82 -861 86 -836
rect 90 -861 94 -836
rect 98 -861 102 -836
rect 120 -861 124 -836
rect 128 -861 132 -836
rect 164 -861 168 -836
rect 172 -861 176 -836
rect 209 -861 213 -836
rect 217 -861 221 -836
rect 329 -907 333 -867
rect 337 -907 341 -867
rect 575 -868 579 -856
rect 584 -868 588 -856
rect 593 -868 597 -856
rect 399 -902 403 -882
rect 407 -902 411 -882
rect 442 -908 446 -868
rect 450 -908 454 -868
rect 615 -869 619 -857
rect 623 -869 627 -857
rect 366 -935 370 -915
rect 374 -935 378 -915
<< polysilicon >>
rect -194 70 -192 73
rect -186 70 -184 73
rect -156 70 -154 73
rect -112 70 -110 73
rect -67 70 -65 73
rect 19 70 21 73
rect 27 70 29 73
rect 57 70 59 73
rect 101 70 103 73
rect 146 70 148 73
rect 512 50 514 53
rect 522 50 524 53
rect -194 38 -192 45
rect -199 34 -192 38
rect -198 23 -196 34
rect -186 26 -184 45
rect -156 37 -154 45
rect -112 37 -110 45
rect -162 35 -154 37
rect -118 35 -110 37
rect -162 23 -160 35
rect -154 23 -152 32
rect -118 23 -116 35
rect -110 23 -108 32
rect -67 23 -65 45
rect 19 38 21 45
rect 14 34 21 38
rect 15 23 17 34
rect 27 26 29 45
rect 57 37 59 45
rect 101 37 103 45
rect 51 35 59 37
rect 95 35 103 37
rect 51 23 53 35
rect 59 23 61 32
rect 95 23 97 35
rect 103 23 105 32
rect 146 23 148 45
rect 266 39 268 43
rect -198 10 -196 13
rect -162 10 -160 13
rect -154 10 -152 13
rect -118 10 -116 13
rect -110 10 -108 13
rect -67 10 -65 13
rect 15 10 17 13
rect 51 10 53 13
rect 59 10 61 13
rect 95 10 97 13
rect 103 10 105 13
rect 146 10 148 13
rect 379 38 381 42
rect 552 49 554 52
rect 303 31 305 38
rect 336 24 338 38
rect 303 8 305 11
rect 336 1 338 4
rect 266 -21 268 -1
rect 512 18 514 38
rect 522 18 524 38
rect 552 23 554 37
rect 552 14 554 17
rect 512 3 514 6
rect 522 3 524 6
rect 303 -9 305 -6
rect 336 -16 338 -13
rect 266 -44 268 -41
rect 303 -43 305 -29
rect 379 -22 381 -2
rect 336 -43 338 -36
rect 379 -45 381 -42
rect -179 -259 -177 -256
rect -171 -259 -169 -256
rect -141 -259 -139 -256
rect -97 -259 -95 -256
rect -52 -259 -50 -256
rect 34 -259 36 -256
rect 42 -259 44 -256
rect 72 -259 74 -256
rect 116 -259 118 -256
rect 161 -259 163 -256
rect 527 -279 529 -276
rect 537 -279 539 -276
rect -179 -291 -177 -284
rect -184 -295 -177 -291
rect -183 -306 -181 -295
rect -171 -303 -169 -284
rect -141 -292 -139 -284
rect -97 -292 -95 -284
rect -147 -294 -139 -292
rect -103 -294 -95 -292
rect -147 -306 -145 -294
rect -139 -306 -137 -297
rect -103 -306 -101 -294
rect -95 -306 -93 -297
rect -52 -306 -50 -284
rect 34 -291 36 -284
rect 29 -295 36 -291
rect 30 -306 32 -295
rect 42 -303 44 -284
rect 72 -292 74 -284
rect 116 -292 118 -284
rect 66 -294 74 -292
rect 110 -294 118 -292
rect 66 -306 68 -294
rect 74 -306 76 -297
rect 110 -306 112 -294
rect 118 -306 120 -297
rect 161 -306 163 -284
rect 281 -290 283 -286
rect -183 -319 -181 -316
rect -147 -319 -145 -316
rect -139 -319 -137 -316
rect -103 -319 -101 -316
rect -95 -319 -93 -316
rect -52 -319 -50 -316
rect 30 -319 32 -316
rect 66 -319 68 -316
rect 74 -319 76 -316
rect 110 -319 112 -316
rect 118 -319 120 -316
rect 161 -319 163 -316
rect 394 -291 396 -287
rect 567 -280 569 -277
rect 318 -298 320 -291
rect 351 -305 353 -291
rect 318 -321 320 -318
rect 351 -328 353 -325
rect 281 -350 283 -330
rect 527 -311 529 -291
rect 537 -311 539 -291
rect 567 -306 569 -292
rect 567 -315 569 -312
rect 527 -326 529 -323
rect 537 -326 539 -323
rect 318 -338 320 -335
rect 351 -345 353 -342
rect 281 -373 283 -370
rect 318 -372 320 -358
rect 394 -351 396 -331
rect 351 -372 353 -365
rect 394 -374 396 -371
rect -155 -526 -153 -523
rect -147 -526 -145 -523
rect -117 -526 -115 -523
rect -73 -526 -71 -523
rect -28 -526 -26 -523
rect 58 -526 60 -523
rect 66 -526 68 -523
rect 96 -526 98 -523
rect 140 -526 142 -523
rect 185 -526 187 -523
rect 551 -546 553 -543
rect 561 -546 563 -543
rect -155 -558 -153 -551
rect -160 -562 -153 -558
rect -159 -573 -157 -562
rect -147 -570 -145 -551
rect -117 -559 -115 -551
rect -73 -559 -71 -551
rect -123 -561 -115 -559
rect -79 -561 -71 -559
rect -123 -573 -121 -561
rect -115 -573 -113 -564
rect -79 -573 -77 -561
rect -71 -573 -69 -564
rect -28 -573 -26 -551
rect 58 -558 60 -551
rect 53 -562 60 -558
rect 54 -573 56 -562
rect 66 -570 68 -551
rect 96 -559 98 -551
rect 140 -559 142 -551
rect 90 -561 98 -559
rect 134 -561 142 -559
rect 90 -573 92 -561
rect 98 -573 100 -564
rect 134 -573 136 -561
rect 142 -573 144 -564
rect 185 -573 187 -551
rect 305 -557 307 -553
rect -159 -586 -157 -583
rect -123 -586 -121 -583
rect -115 -586 -113 -583
rect -79 -586 -77 -583
rect -71 -586 -69 -583
rect -28 -586 -26 -583
rect 54 -586 56 -583
rect 90 -586 92 -583
rect 98 -586 100 -583
rect 134 -586 136 -583
rect 142 -586 144 -583
rect 185 -586 187 -583
rect 418 -558 420 -554
rect 591 -547 593 -544
rect 342 -565 344 -558
rect 375 -572 377 -558
rect 342 -588 344 -585
rect 375 -595 377 -592
rect 305 -617 307 -597
rect 551 -578 553 -558
rect 561 -578 563 -558
rect 591 -573 593 -559
rect 591 -582 593 -579
rect 551 -593 553 -590
rect 561 -593 563 -590
rect 342 -605 344 -602
rect 375 -612 377 -609
rect 305 -640 307 -637
rect 342 -639 344 -625
rect 418 -618 420 -598
rect 375 -639 377 -632
rect 418 -641 420 -638
rect -126 -836 -124 -833
rect -118 -836 -116 -833
rect -88 -836 -86 -833
rect -44 -836 -42 -833
rect 1 -836 3 -833
rect 87 -836 89 -833
rect 95 -836 97 -833
rect 125 -836 127 -833
rect 169 -836 171 -833
rect 214 -836 216 -833
rect 580 -856 582 -853
rect 590 -856 592 -853
rect -126 -868 -124 -861
rect -131 -872 -124 -868
rect -130 -883 -128 -872
rect -118 -880 -116 -861
rect -88 -869 -86 -861
rect -44 -869 -42 -861
rect -94 -871 -86 -869
rect -50 -871 -42 -869
rect -94 -883 -92 -871
rect -86 -883 -84 -874
rect -50 -883 -48 -871
rect -42 -883 -40 -874
rect 1 -883 3 -861
rect 87 -868 89 -861
rect 82 -872 89 -868
rect 83 -883 85 -872
rect 95 -880 97 -861
rect 125 -869 127 -861
rect 169 -869 171 -861
rect 119 -871 127 -869
rect 163 -871 171 -869
rect 119 -883 121 -871
rect 127 -883 129 -874
rect 163 -883 165 -871
rect 171 -883 173 -874
rect 214 -883 216 -861
rect 334 -867 336 -863
rect -130 -896 -128 -893
rect -94 -896 -92 -893
rect -86 -896 -84 -893
rect -50 -896 -48 -893
rect -42 -896 -40 -893
rect 1 -896 3 -893
rect 83 -896 85 -893
rect 119 -896 121 -893
rect 127 -896 129 -893
rect 163 -896 165 -893
rect 171 -896 173 -893
rect 214 -896 216 -893
rect 447 -868 449 -864
rect 620 -857 622 -854
rect 371 -875 373 -868
rect 404 -882 406 -868
rect 371 -898 373 -895
rect 404 -905 406 -902
rect 334 -927 336 -907
rect 580 -888 582 -868
rect 590 -888 592 -868
rect 620 -883 622 -869
rect 620 -892 622 -889
rect 580 -903 582 -900
rect 590 -903 592 -900
rect 371 -915 373 -912
rect 404 -922 406 -919
rect 334 -950 336 -947
rect 371 -949 373 -935
rect 447 -928 449 -908
rect 404 -949 406 -942
rect 447 -951 449 -948
<< polycontact >>
rect -203 34 -199 38
rect -190 26 -186 30
rect -167 26 -162 31
rect -152 26 -147 30
rect -123 26 -118 31
rect -71 31 -67 36
rect -108 26 -103 30
rect 10 34 14 38
rect 23 26 27 30
rect 46 26 51 31
rect 61 26 66 30
rect 90 26 95 31
rect 142 31 146 36
rect 105 26 110 30
rect 302 38 306 43
rect 335 38 339 43
rect 262 -18 266 -13
rect 508 27 512 31
rect 518 21 522 25
rect 548 26 552 30
rect 375 -19 379 -14
rect 302 -48 306 -43
rect 335 -48 339 -43
rect -188 -295 -184 -291
rect -175 -303 -171 -299
rect -152 -303 -147 -298
rect -137 -303 -132 -299
rect -108 -303 -103 -298
rect -56 -298 -52 -293
rect -93 -303 -88 -299
rect 25 -295 29 -291
rect 38 -303 42 -299
rect 61 -303 66 -298
rect 76 -303 81 -299
rect 105 -303 110 -298
rect 157 -298 161 -293
rect 120 -303 125 -299
rect 317 -291 321 -286
rect 350 -291 354 -286
rect 277 -347 281 -342
rect 523 -302 527 -298
rect 533 -308 537 -304
rect 563 -303 567 -299
rect 390 -348 394 -343
rect 317 -377 321 -372
rect 350 -377 354 -372
rect -164 -562 -160 -558
rect -151 -570 -147 -566
rect -128 -570 -123 -565
rect -113 -570 -108 -566
rect -84 -570 -79 -565
rect -32 -565 -28 -560
rect -69 -570 -64 -566
rect 49 -562 53 -558
rect 62 -570 66 -566
rect 85 -570 90 -565
rect 100 -570 105 -566
rect 129 -570 134 -565
rect 181 -565 185 -560
rect 144 -570 149 -566
rect 341 -558 345 -553
rect 374 -558 378 -553
rect 301 -614 305 -609
rect 547 -569 551 -565
rect 557 -575 561 -571
rect 587 -570 591 -566
rect 414 -615 418 -610
rect 341 -644 345 -639
rect 374 -644 378 -639
rect -135 -872 -131 -868
rect -122 -880 -118 -876
rect -99 -880 -94 -875
rect -84 -880 -79 -876
rect -55 -880 -50 -875
rect -3 -875 1 -870
rect -40 -880 -35 -876
rect 78 -872 82 -868
rect 91 -880 95 -876
rect 114 -880 119 -875
rect 129 -880 134 -876
rect 158 -880 163 -875
rect 210 -875 214 -870
rect 173 -880 178 -876
rect 370 -868 374 -863
rect 403 -868 407 -863
rect 330 -924 334 -919
rect 576 -879 580 -875
rect 586 -885 590 -881
rect 616 -880 620 -876
rect 443 -925 447 -920
rect 370 -954 374 -949
rect 403 -954 407 -949
<< metal1 >>
rect -205 76 499 80
rect -199 70 -195 76
rect -161 70 -157 76
rect -117 70 -113 76
rect -72 70 -68 76
rect 14 70 18 76
rect 52 70 56 76
rect 96 70 100 76
rect 141 70 145 76
rect 233 75 499 76
rect -149 45 -136 70
rect -105 45 -92 70
rect 64 45 77 70
rect 108 45 121 70
rect -210 34 -203 38
rect -183 37 -179 45
rect -183 34 -143 37
rect -193 26 -190 30
rect -183 23 -179 34
rect -171 26 -167 31
rect -147 26 -143 34
rect -139 31 -136 45
rect -95 36 -92 45
rect -95 31 -71 36
rect -64 35 -60 45
rect -139 26 -123 31
rect -103 26 -99 30
rect -139 23 -136 26
rect -95 23 -92 31
rect -64 30 -51 35
rect -64 23 -60 30
rect 3 34 10 38
rect 30 37 34 45
rect 30 34 70 37
rect 20 26 23 30
rect 30 23 34 34
rect 42 26 46 31
rect 66 26 70 34
rect 74 31 77 45
rect 118 36 121 45
rect 118 31 142 36
rect 149 35 153 45
rect 261 39 265 75
rect 74 26 90 31
rect 110 26 114 30
rect 74 23 77 26
rect 118 23 121 31
rect 149 30 162 35
rect 149 23 153 30
rect -191 13 -179 23
rect -147 13 -136 23
rect -103 13 -92 23
rect 22 13 34 23
rect 66 13 77 23
rect 110 13 121 23
rect -203 8 -199 13
rect -167 8 -163 13
rect -123 8 -119 13
rect -72 8 -68 13
rect 10 8 14 13
rect 46 8 50 13
rect 90 8 94 13
rect 141 8 145 13
rect -204 4 153 8
rect 149 -81 153 4
rect 286 7 291 62
rect 302 43 306 50
rect 335 43 339 50
rect 374 38 378 75
rect 461 55 467 62
rect 494 59 499 75
rect 494 58 544 59
rect 494 56 565 58
rect 394 50 475 55
rect 298 7 302 11
rect 286 3 302 7
rect 252 -18 262 -13
rect 269 -14 273 -1
rect 298 -9 302 3
rect 269 -19 282 -14
rect 269 -21 273 -19
rect 306 6 310 11
rect 306 2 323 6
rect 306 -9 310 2
rect 319 -8 323 2
rect 331 -8 335 4
rect 319 -13 335 -8
rect 261 -80 265 -41
rect 302 -61 306 -48
rect 319 -74 325 -13
rect 331 -16 335 -13
rect 339 -9 343 4
rect 339 -13 360 -9
rect 339 -16 343 -13
rect 354 -14 360 -13
rect 354 -19 364 -14
rect 370 -19 375 -14
rect 382 -15 386 -2
rect 424 24 433 37
rect 472 30 475 50
rect 507 50 510 56
rect 526 50 529 56
rect 541 55 565 56
rect 547 49 550 55
rect 516 35 519 38
rect 516 32 529 35
rect 472 27 508 30
rect 526 29 529 32
rect 526 26 548 29
rect 556 29 559 37
rect 556 26 568 29
rect 424 21 518 24
rect 382 -20 399 -15
rect 382 -22 386 -20
rect 335 -61 339 -48
rect 374 -80 378 -42
rect 424 -60 432 21
rect 526 18 529 26
rect 556 23 559 26
rect 547 13 550 17
rect 537 10 565 13
rect 507 0 510 6
rect 537 0 541 10
rect 442 -3 541 0
rect 442 -80 453 -3
rect 233 -81 453 -80
rect 149 -88 453 -81
rect -190 -253 514 -249
rect -184 -259 -180 -253
rect -146 -259 -142 -253
rect -102 -259 -98 -253
rect -57 -259 -53 -253
rect 29 -259 33 -253
rect 67 -259 71 -253
rect 111 -259 115 -253
rect 156 -259 160 -253
rect 248 -254 514 -253
rect -134 -284 -121 -259
rect -90 -284 -77 -259
rect 79 -284 92 -259
rect 123 -284 136 -259
rect -195 -295 -188 -291
rect -168 -292 -164 -284
rect -168 -295 -128 -292
rect -178 -303 -175 -299
rect -168 -306 -164 -295
rect -156 -303 -152 -298
rect -132 -303 -128 -295
rect -124 -298 -121 -284
rect -80 -293 -77 -284
rect -80 -298 -56 -293
rect -49 -294 -45 -284
rect -124 -303 -108 -298
rect -88 -303 -84 -299
rect -124 -306 -121 -303
rect -80 -306 -77 -298
rect -49 -299 -36 -294
rect -49 -306 -45 -299
rect 18 -295 25 -291
rect 45 -292 49 -284
rect 45 -295 85 -292
rect 35 -303 38 -299
rect 45 -306 49 -295
rect 57 -303 61 -298
rect 81 -303 85 -295
rect 89 -298 92 -284
rect 133 -293 136 -284
rect 133 -298 157 -293
rect 164 -294 168 -284
rect 276 -290 280 -254
rect 89 -303 105 -298
rect 125 -303 129 -299
rect 89 -306 92 -303
rect 133 -306 136 -298
rect 164 -299 177 -294
rect 164 -306 168 -299
rect -176 -316 -164 -306
rect -132 -316 -121 -306
rect -88 -316 -77 -306
rect 37 -316 49 -306
rect 81 -316 92 -306
rect 125 -316 136 -306
rect -188 -321 -184 -316
rect -152 -321 -148 -316
rect -108 -321 -104 -316
rect -57 -321 -53 -316
rect 25 -321 29 -316
rect 61 -321 65 -316
rect 105 -321 109 -316
rect 156 -321 160 -316
rect -189 -325 168 -321
rect 164 -410 168 -325
rect 301 -322 306 -267
rect 317 -286 321 -279
rect 350 -286 354 -279
rect 389 -291 393 -254
rect 476 -274 482 -267
rect 509 -270 514 -254
rect 509 -271 559 -270
rect 509 -273 580 -271
rect 409 -279 490 -274
rect 313 -322 317 -318
rect 301 -326 317 -322
rect 267 -347 277 -342
rect 284 -343 288 -330
rect 313 -338 317 -326
rect 284 -348 297 -343
rect 284 -350 288 -348
rect 321 -323 325 -318
rect 321 -327 338 -323
rect 321 -338 325 -327
rect 334 -337 338 -327
rect 346 -337 350 -325
rect 334 -342 350 -337
rect 276 -409 280 -370
rect 317 -390 321 -377
rect 334 -403 340 -342
rect 346 -345 350 -342
rect 354 -338 358 -325
rect 354 -342 375 -338
rect 354 -345 358 -342
rect 369 -343 375 -342
rect 369 -348 379 -343
rect 385 -348 390 -343
rect 397 -344 401 -331
rect 439 -305 448 -292
rect 487 -299 490 -279
rect 522 -279 525 -273
rect 541 -279 544 -273
rect 556 -274 580 -273
rect 562 -280 565 -274
rect 531 -294 534 -291
rect 531 -297 544 -294
rect 487 -302 523 -299
rect 541 -300 544 -297
rect 541 -303 563 -300
rect 571 -300 574 -292
rect 571 -303 583 -300
rect 439 -308 533 -305
rect 397 -349 414 -344
rect 397 -351 401 -349
rect 350 -390 354 -377
rect 389 -409 393 -371
rect 439 -389 447 -308
rect 541 -311 544 -303
rect 571 -306 574 -303
rect 562 -316 565 -312
rect 552 -319 580 -316
rect 522 -329 525 -323
rect 552 -329 556 -319
rect 457 -332 556 -329
rect 457 -409 468 -332
rect 248 -410 468 -409
rect 164 -417 468 -410
rect -166 -520 538 -516
rect -160 -526 -156 -520
rect -122 -526 -118 -520
rect -78 -526 -74 -520
rect -33 -526 -29 -520
rect 53 -526 57 -520
rect 91 -526 95 -520
rect 135 -526 139 -520
rect 180 -526 184 -520
rect 272 -521 538 -520
rect -110 -551 -97 -526
rect -66 -551 -53 -526
rect 103 -551 116 -526
rect 147 -551 160 -526
rect -171 -562 -164 -558
rect -144 -559 -140 -551
rect -144 -562 -104 -559
rect -154 -570 -151 -566
rect -144 -573 -140 -562
rect -132 -570 -128 -565
rect -108 -570 -104 -562
rect -100 -565 -97 -551
rect -56 -560 -53 -551
rect -56 -565 -32 -560
rect -25 -561 -21 -551
rect -100 -570 -84 -565
rect -64 -570 -60 -566
rect -100 -573 -97 -570
rect -56 -573 -53 -565
rect -25 -566 -12 -561
rect -25 -573 -21 -566
rect 42 -562 49 -558
rect 69 -559 73 -551
rect 69 -562 109 -559
rect 59 -570 62 -566
rect 69 -573 73 -562
rect 81 -570 85 -565
rect 105 -570 109 -562
rect 113 -565 116 -551
rect 157 -560 160 -551
rect 157 -565 181 -560
rect 188 -561 192 -551
rect 300 -557 304 -521
rect 113 -570 129 -565
rect 149 -570 153 -566
rect 113 -573 116 -570
rect 157 -573 160 -565
rect 188 -566 201 -561
rect 188 -573 192 -566
rect -152 -583 -140 -573
rect -108 -583 -97 -573
rect -64 -583 -53 -573
rect 61 -583 73 -573
rect 105 -583 116 -573
rect 149 -583 160 -573
rect -164 -588 -160 -583
rect -128 -588 -124 -583
rect -84 -588 -80 -583
rect -33 -588 -29 -583
rect 49 -588 53 -583
rect 85 -588 89 -583
rect 129 -588 133 -583
rect 180 -588 184 -583
rect -165 -592 192 -588
rect 188 -677 192 -592
rect 325 -589 330 -534
rect 341 -553 345 -546
rect 374 -553 378 -546
rect 413 -558 417 -521
rect 500 -541 506 -534
rect 533 -537 538 -521
rect 533 -538 583 -537
rect 533 -540 604 -538
rect 433 -546 514 -541
rect 337 -589 341 -585
rect 325 -593 341 -589
rect 291 -614 301 -609
rect 308 -610 312 -597
rect 337 -605 341 -593
rect 308 -615 321 -610
rect 308 -617 312 -615
rect 345 -590 349 -585
rect 345 -594 362 -590
rect 345 -605 349 -594
rect 358 -604 362 -594
rect 370 -604 374 -592
rect 358 -609 374 -604
rect 300 -676 304 -637
rect 341 -657 345 -644
rect 358 -670 364 -609
rect 370 -612 374 -609
rect 378 -605 382 -592
rect 378 -609 399 -605
rect 378 -612 382 -609
rect 393 -610 399 -609
rect 393 -615 403 -610
rect 409 -615 414 -610
rect 421 -611 425 -598
rect 463 -572 472 -559
rect 511 -566 514 -546
rect 546 -546 549 -540
rect 565 -546 568 -540
rect 580 -541 604 -540
rect 586 -547 589 -541
rect 555 -561 558 -558
rect 555 -564 568 -561
rect 511 -569 547 -566
rect 565 -567 568 -564
rect 565 -570 587 -567
rect 595 -567 598 -559
rect 595 -570 607 -567
rect 463 -575 557 -572
rect 421 -616 438 -611
rect 421 -618 425 -616
rect 374 -657 378 -644
rect 413 -676 417 -638
rect 463 -656 471 -575
rect 565 -578 568 -570
rect 595 -573 598 -570
rect 586 -583 589 -579
rect 576 -586 604 -583
rect 546 -596 549 -590
rect 576 -596 580 -586
rect 481 -599 580 -596
rect 481 -676 492 -599
rect 272 -677 492 -676
rect 188 -684 492 -677
rect -137 -830 567 -826
rect -131 -836 -127 -830
rect -93 -836 -89 -830
rect -49 -836 -45 -830
rect -4 -836 0 -830
rect 82 -836 86 -830
rect 120 -836 124 -830
rect 164 -836 168 -830
rect 209 -836 213 -830
rect 301 -831 567 -830
rect -81 -861 -68 -836
rect -37 -861 -24 -836
rect 132 -861 145 -836
rect 176 -861 189 -836
rect -142 -872 -135 -868
rect -115 -869 -111 -861
rect -115 -872 -75 -869
rect -125 -880 -122 -876
rect -115 -883 -111 -872
rect -103 -880 -99 -875
rect -79 -880 -75 -872
rect -71 -875 -68 -861
rect -27 -870 -24 -861
rect -27 -875 -3 -870
rect 4 -871 8 -861
rect -71 -880 -55 -875
rect -35 -880 -31 -876
rect -71 -883 -68 -880
rect -27 -883 -24 -875
rect 4 -876 17 -871
rect 4 -883 8 -876
rect 71 -872 78 -868
rect 98 -869 102 -861
rect 98 -872 138 -869
rect 88 -880 91 -876
rect 98 -883 102 -872
rect 110 -880 114 -875
rect 134 -880 138 -872
rect 142 -875 145 -861
rect 186 -870 189 -861
rect 186 -875 210 -870
rect 217 -871 221 -861
rect 329 -867 333 -831
rect 142 -880 158 -875
rect 178 -880 182 -876
rect 142 -883 145 -880
rect 186 -883 189 -875
rect 217 -876 230 -871
rect 217 -883 221 -876
rect -123 -893 -111 -883
rect -79 -893 -68 -883
rect -35 -893 -24 -883
rect 90 -893 102 -883
rect 134 -893 145 -883
rect 178 -893 189 -883
rect -135 -898 -131 -893
rect -99 -898 -95 -893
rect -55 -898 -51 -893
rect -4 -898 0 -893
rect 78 -898 82 -893
rect 114 -898 118 -893
rect 158 -898 162 -893
rect 209 -898 213 -893
rect -136 -902 221 -898
rect 217 -987 221 -902
rect 354 -899 359 -844
rect 370 -863 374 -856
rect 403 -863 407 -856
rect 442 -868 446 -831
rect 529 -851 535 -844
rect 562 -847 567 -831
rect 562 -848 612 -847
rect 562 -850 633 -848
rect 462 -856 543 -851
rect 366 -899 370 -895
rect 354 -903 370 -899
rect 320 -924 330 -919
rect 337 -920 341 -907
rect 366 -915 370 -903
rect 337 -925 350 -920
rect 337 -927 341 -925
rect 374 -900 378 -895
rect 374 -904 391 -900
rect 374 -915 378 -904
rect 387 -914 391 -904
rect 399 -914 403 -902
rect 387 -919 403 -914
rect 329 -986 333 -947
rect 370 -967 374 -954
rect 387 -980 393 -919
rect 399 -922 403 -919
rect 407 -915 411 -902
rect 407 -919 428 -915
rect 407 -922 411 -919
rect 422 -920 428 -919
rect 422 -925 432 -920
rect 438 -925 443 -920
rect 450 -921 454 -908
rect 492 -882 501 -869
rect 540 -876 543 -856
rect 575 -856 578 -850
rect 594 -856 597 -850
rect 609 -851 633 -850
rect 615 -857 618 -851
rect 584 -871 587 -868
rect 584 -874 597 -871
rect 540 -879 576 -876
rect 594 -877 597 -874
rect 594 -880 616 -877
rect 624 -877 627 -869
rect 624 -880 636 -877
rect 492 -885 586 -882
rect 450 -926 467 -921
rect 450 -928 454 -926
rect 403 -967 407 -954
rect 442 -986 446 -948
rect 492 -966 500 -885
rect 594 -888 597 -880
rect 624 -883 627 -880
rect 615 -893 618 -889
rect 605 -896 633 -893
rect 575 -906 578 -900
rect 605 -906 609 -896
rect 510 -909 609 -906
rect 510 -986 521 -909
rect 301 -987 521 -986
rect 217 -994 521 -987
<< m2contact >>
rect -51 29 -40 36
rect 286 62 292 67
rect 162 29 173 36
rect 302 50 307 55
rect 334 50 339 55
rect 458 62 468 69
rect 386 50 394 55
rect 247 -18 252 -13
rect 282 -19 288 -14
rect 302 -66 307 -61
rect 423 37 434 43
rect 364 -19 370 -14
rect 399 -20 405 -15
rect 335 -66 340 -61
rect 424 -66 432 -60
rect -36 -300 -25 -293
rect 301 -267 307 -262
rect 177 -300 188 -293
rect 317 -279 322 -274
rect 349 -279 354 -274
rect 473 -267 483 -260
rect 401 -279 409 -274
rect 262 -347 267 -342
rect 297 -348 303 -343
rect 317 -395 322 -390
rect 438 -292 449 -286
rect 379 -348 385 -343
rect 414 -349 420 -344
rect 350 -395 355 -390
rect 439 -395 447 -389
rect -12 -567 -1 -560
rect 325 -534 331 -529
rect 201 -567 212 -560
rect 341 -546 346 -541
rect 373 -546 378 -541
rect 497 -534 507 -527
rect 425 -546 433 -541
rect 286 -614 291 -609
rect 321 -615 327 -610
rect 341 -662 346 -657
rect 462 -559 473 -553
rect 403 -615 409 -610
rect 438 -616 444 -611
rect 374 -662 379 -657
rect 463 -662 471 -656
rect 17 -877 28 -870
rect 354 -844 360 -839
rect 230 -877 241 -870
rect 370 -856 375 -851
rect 402 -856 407 -851
rect 526 -844 536 -837
rect 454 -856 462 -851
rect 315 -924 320 -919
rect 350 -925 356 -920
rect 370 -972 375 -967
rect 491 -869 502 -863
rect 432 -925 438 -920
rect 467 -926 473 -921
rect 403 -972 408 -967
rect 492 -972 500 -966
<< metal2 >>
rect 188 98 192 99
rect 188 94 466 98
rect -25 83 170 87
rect -25 35 -21 83
rect -40 30 -21 35
rect 188 35 192 94
rect 231 85 431 89
rect 292 62 405 67
rect 173 30 192 35
rect 247 50 302 55
rect 307 50 334 55
rect 339 50 386 55
rect 247 -13 251 50
rect 282 -61 288 -19
rect 364 -60 370 -19
rect 399 -15 405 62
rect 425 43 431 85
rect 461 69 466 94
rect 281 -66 302 -61
rect 307 -66 335 -61
rect 340 -66 354 -61
rect 364 -66 424 -60
rect 203 -231 207 -230
rect 203 -235 481 -231
rect -10 -246 185 -242
rect -10 -294 -6 -246
rect -25 -299 -6 -294
rect 203 -294 207 -235
rect 246 -244 446 -240
rect 307 -267 420 -262
rect 188 -299 207 -294
rect 262 -279 317 -274
rect 322 -279 349 -274
rect 354 -279 401 -274
rect 262 -342 266 -279
rect 297 -390 303 -348
rect 379 -389 385 -348
rect 414 -344 420 -267
rect 440 -286 446 -244
rect 476 -260 481 -235
rect 296 -395 317 -390
rect 322 -395 350 -390
rect 355 -395 369 -390
rect 379 -395 439 -389
rect 227 -498 231 -497
rect 227 -502 505 -498
rect 14 -513 209 -509
rect 14 -561 18 -513
rect -1 -566 18 -561
rect 227 -561 231 -502
rect 270 -511 470 -507
rect 331 -534 444 -529
rect 212 -566 231 -561
rect 286 -546 341 -541
rect 346 -546 373 -541
rect 378 -546 425 -541
rect 286 -609 290 -546
rect 321 -657 327 -615
rect 403 -656 409 -615
rect 438 -611 444 -534
rect 464 -553 470 -511
rect 500 -527 505 -502
rect 320 -662 341 -657
rect 346 -662 374 -657
rect 379 -662 393 -657
rect 403 -662 463 -656
rect 256 -808 260 -807
rect 256 -812 534 -808
rect 43 -823 238 -819
rect 43 -871 47 -823
rect 28 -876 47 -871
rect 256 -871 260 -812
rect 299 -821 499 -817
rect 360 -844 473 -839
rect 241 -876 260 -871
rect 315 -856 370 -851
rect 375 -856 402 -851
rect 407 -856 454 -851
rect 315 -919 319 -856
rect 350 -967 356 -925
rect 432 -966 438 -925
rect 467 -921 473 -844
rect 493 -863 499 -821
rect 529 -837 534 -812
rect 349 -972 370 -967
rect 375 -972 403 -967
rect 408 -972 422 -967
rect 432 -972 492 -966
<< m3contact >>
rect 170 82 183 88
rect 221 83 231 89
rect 185 -247 198 -241
rect 236 -246 246 -240
rect 209 -514 222 -508
rect 260 -513 270 -507
rect 238 -824 251 -818
rect 289 -823 299 -817
<< metal3 >>
rect 183 83 221 88
rect 198 -246 236 -241
rect 222 -513 260 -508
rect 251 -823 289 -818
<< labels >>
rlabel metal1 563 26 568 29 1 g0
rlabel metal1 501 21 504 24 1 b0_reg
rlabel metal1 501 27 505 30 1 a0_reg
rlabel metal1 561 11 561 11 1 gnd!
rlabel metal1 555 56 555 56 5 vdd!
rlabel metal1 525 -2 525 -2 1 gnd!
rlabel metal1 525 58 525 58 5 vdd!
rlabel metal1 458 50 473 55 1 a0_reg
rlabel metal1 424 -1 432 15 1 b0_reg
rlabel metal1 319 -73 325 -67 1 p0
rlabel metal1 342 75 456 80 1 vdd
rlabel metal1 318 -87 432 -81 1 gnd
rlabel metal1 20 27 22 29 1 clk
rlabel metal1 18 6 21 7 1 gnd
rlabel metal1 24 78 26 79 5 vdd
rlabel metal1 43 27 44 29 1 clk
rlabel metal1 111 27 113 29 1 clk
rlabel metal1 155 32 158 34 1 a0_reg
rlabel metal1 5 35 7 37 3 a0
rlabel metal1 -102 27 -100 29 1 clk
rlabel metal1 -170 27 -169 29 1 clk
rlabel metal1 -189 78 -187 79 5 vdd
rlabel metal1 -195 6 -192 7 1 gnd
rlabel metal1 -193 27 -191 29 1 clk
rlabel metal1 -208 35 -206 37 3 b0
rlabel metal1 -58 32 -55 34 1 b0_reg
rlabel metal1 576 -318 576 -318 1 gnd!
rlabel metal1 570 -273 570 -273 5 vdd!
rlabel metal1 540 -331 540 -331 1 gnd!
rlabel metal1 540 -271 540 -271 5 vdd!
rlabel metal1 357 -254 471 -249 1 vdd
rlabel metal1 333 -416 447 -410 1 gnd
rlabel metal1 35 -302 37 -300 1 clk
rlabel metal1 33 -323 36 -322 1 gnd
rlabel metal1 39 -251 41 -250 5 vdd
rlabel metal1 58 -302 59 -300 1 clk
rlabel metal1 126 -302 128 -300 1 clk
rlabel metal1 -87 -302 -85 -300 1 clk
rlabel metal1 -155 -302 -154 -300 1 clk
rlabel metal1 -174 -251 -172 -250 5 vdd
rlabel metal1 -180 -323 -177 -322 1 gnd
rlabel metal1 -178 -302 -176 -300 1 clk
rlabel metal1 600 -585 600 -585 1 gnd!
rlabel metal1 594 -540 594 -540 5 vdd!
rlabel metal1 564 -598 564 -598 1 gnd!
rlabel metal1 564 -538 564 -538 5 vdd!
rlabel metal1 381 -521 495 -516 1 vdd
rlabel metal1 357 -683 471 -677 1 gnd
rlabel metal1 59 -569 61 -567 1 clk
rlabel metal1 57 -590 60 -589 1 gnd
rlabel metal1 63 -518 65 -517 5 vdd
rlabel metal1 82 -569 83 -567 1 clk
rlabel metal1 150 -569 152 -567 1 clk
rlabel metal1 -63 -569 -61 -567 1 clk
rlabel metal1 -131 -569 -130 -567 1 clk
rlabel metal1 -150 -518 -148 -517 5 vdd
rlabel metal1 -156 -590 -153 -589 1 gnd
rlabel metal1 -154 -569 -152 -567 1 clk
rlabel metal1 -125 -879 -123 -877 1 clk
rlabel metal1 -127 -900 -124 -899 1 gnd
rlabel metal1 -121 -828 -119 -827 5 vdd
rlabel metal1 -102 -879 -101 -877 1 clk
rlabel metal1 -34 -879 -32 -877 1 clk
rlabel metal1 179 -879 181 -877 1 clk
rlabel metal1 111 -879 112 -877 1 clk
rlabel metal1 92 -828 94 -827 5 vdd
rlabel metal1 86 -900 89 -899 1 gnd
rlabel metal1 88 -879 90 -877 1 clk
rlabel metal1 386 -993 500 -987 1 gnd
rlabel metal1 410 -831 524 -826 1 vdd
rlabel metal1 593 -848 593 -848 5 vdd!
rlabel metal1 593 -908 593 -908 1 gnd!
rlabel metal1 623 -850 623 -850 5 vdd!
rlabel metal1 629 -895 629 -895 1 gnd!
rlabel metal1 20 -294 22 -292 1 a1
rlabel metal1 -45 -297 -40 -295 1 b1_reg
rlabel metal1 -193 -294 -191 -292 1 b1
rlabel metal1 170 -297 173 -295 1 a1_reg
rlabel metal1 334 -402 340 -396 1 p1
rlabel metal1 473 -279 488 -274 1 a1_reg
rlabel metal1 516 -308 519 -305 1 b1_reg
rlabel metal1 516 -302 520 -299 1 a1_reg
rlabel metal1 578 -303 583 -300 1 g1
rlabel metal1 44 -561 46 -559 1 a2
rlabel metal1 194 -564 197 -562 1 a2_reg
rlabel metal1 -19 -564 -16 -562 1 b2_reg
rlabel metal1 -169 -561 -166 -559 1 b2
rlabel metal1 497 -546 512 -541 1 a2_reg
rlabel metal1 540 -569 544 -566 1 a2_reg
rlabel metal1 540 -575 544 -572 1 b2_reg
rlabel metal1 358 -669 364 -663 1 p2
rlabel metal1 602 -570 607 -567 1 g2
rlabel metal1 631 -880 636 -877 7 g3
rlabel metal1 569 -879 574 -876 1 a3_reg
rlabel metal1 569 -885 574 -882 1 b3_reg
rlabel metal1 463 -597 471 -581 1 b2_reg
rlabel metal1 439 -330 447 -313 1 b1_reg
rlabel metal1 492 -908 500 -891 1 b3_reg
rlabel metal1 526 -856 541 -851 1 a3_reg
rlabel metal1 387 -979 393 -973 1 p3
rlabel metal1 223 -874 226 -872 1 a3_reg
rlabel metal1 73 -871 76 -869 1 a3
rlabel metal1 10 -874 13 -872 1 b3_reg
rlabel metal1 -140 -871 -137 -869 1 b3
<< end >>
