.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd
.option scale=0.09u
Vdd    vdd gnd 'SUPPLY'
vin    a 0 pulse 0 1.8 0ns 0ns 0ns 15ns 30ns  
vin2   b 0 pulse 0 1.8 0ns 0ns 0ns 24ns 48ns 

M1000 a_13_n26# a gnd Gnd CMOSN w=12 l=2
+  ad=96 pd=40 as=90 ps=56
M1001 in a vdd w_0_0# CMOSP w=12 l=2
+  ad=96 pd=40 as=180 ps=102
M1002 op in vdd w_40_n1# CMOSP w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1003 vdd b in w_0_0# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 op in gnd Gnd CMOSN w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1005 in b a_13_n26# Gnd CMOSN w=12 l=2
+  ad=60 pd=34 as=0 ps=0
C0 a w_0_0# 0.06fF
C1 w_0_0# in 0.04fF
C2 gnd op 0.10fF
C3 gnd in 0.08fF
C4 op in 0.04fF
C5 w_40_n1# op 0.03fF
C6 w_40_n1# in 0.06fF
C7 w_0_0# b 0.06fF
C8 a b 0.24fF
C9 gnd b 0.05fF
C10 in b 0.13fF
C11 vdd w_0_0# 0.10fF
C12 vdd a 0.02fF
C13 vdd op 0.15fF
C14 vdd in 0.30fF
C15 w_40_n1# vdd 0.06fF
C16 gnd Gnd 0.27fF
C17 op Gnd 0.05fF
C18 in Gnd 0.23fF
C19 vdd Gnd 0.12fF
C20 b Gnd 0.20fF
C21 a Gnd 0.17fF
C22 w_40_n1# Gnd 0.58fF
C23 w_0_0# Gnd 0.82fF


    .tran 0.1n 200n
    .control
    run
     set curplottitle  = "Eswar-2023102011"
    plot 5+v(a) 3+v(b) v(op)
    .endc
