magic
tech scmos
timestamp 1731734105
<< nwell >>
rect -206 21 -174 58
rect -168 21 -142 58
rect -124 21 -98 58
rect -79 21 -53 58
rect 7 21 39 58
rect 45 21 71 58
rect 89 21 115 58
rect 134 21 160 58
rect 254 -29 279 28
rect 291 -57 316 -17
rect 324 -24 349 16
rect 367 -30 392 27
rect 500 14 534 38
rect 540 13 564 37
<< ntransistor >>
rect -199 -5 -197 5
rect -163 -5 -161 5
rect -155 -5 -153 5
rect -119 -5 -117 5
rect -111 -5 -109 5
rect -68 -5 -66 5
rect 14 -5 16 5
rect 50 -5 52 5
rect 58 -5 60 5
rect 94 -5 96 5
rect 102 -5 104 5
rect 145 -5 147 5
rect 302 -7 304 13
rect 511 -12 513 0
rect 521 -12 523 0
rect 551 -1 553 5
rect 265 -59 267 -39
rect 335 -54 337 -34
rect 378 -60 380 -40
<< ptransistor >>
rect -195 27 -193 52
rect -187 27 -185 52
rect -157 27 -155 52
rect -113 27 -111 52
rect -68 27 -66 52
rect 18 27 20 52
rect 26 27 28 52
rect 56 27 58 52
rect 100 27 102 52
rect 145 27 147 52
rect 265 -19 267 21
rect 511 20 513 32
rect 521 20 523 32
rect 335 -14 337 6
rect 378 -20 380 20
rect 551 19 553 31
rect 302 -47 304 -27
<< ndiffusion >>
rect -200 -5 -199 5
rect -197 -5 -196 5
rect -164 -5 -163 5
rect -161 -5 -160 5
rect -156 -5 -155 5
rect -153 -5 -152 5
rect -120 -5 -119 5
rect -117 -5 -116 5
rect -112 -5 -111 5
rect -109 -5 -108 5
rect -69 -5 -68 5
rect -66 -5 -65 5
rect 13 -5 14 5
rect 16 -5 17 5
rect 49 -5 50 5
rect 52 -5 53 5
rect 57 -5 58 5
rect 60 -5 61 5
rect 93 -5 94 5
rect 96 -5 97 5
rect 101 -5 102 5
rect 104 -5 105 5
rect 144 -5 145 5
rect 147 -5 148 5
rect 301 -7 302 13
rect 304 -7 305 13
rect 510 -12 511 0
rect 513 -12 521 0
rect 523 -12 524 0
rect 550 -1 551 5
rect 553 -1 554 5
rect 264 -59 265 -39
rect 267 -59 268 -39
rect 334 -54 335 -34
rect 337 -54 338 -34
rect 377 -60 378 -40
rect 380 -60 381 -40
<< pdiffusion >>
rect -196 27 -195 52
rect -193 27 -192 52
rect -188 27 -187 52
rect -185 27 -184 52
rect -158 27 -157 52
rect -155 27 -154 52
rect -114 27 -113 52
rect -111 27 -110 52
rect -69 27 -68 52
rect -66 27 -65 52
rect 17 27 18 52
rect 20 27 21 52
rect 25 27 26 52
rect 28 27 29 52
rect 55 27 56 52
rect 58 27 59 52
rect 99 27 100 52
rect 102 27 103 52
rect 144 27 145 52
rect 147 27 148 52
rect 264 -19 265 21
rect 267 -19 268 21
rect 510 20 511 32
rect 513 20 515 32
rect 519 20 521 32
rect 523 20 524 32
rect 334 -14 335 6
rect 337 -14 338 6
rect 377 -20 378 20
rect 380 -20 381 20
rect 550 19 551 31
rect 553 19 554 31
rect 301 -47 302 -27
rect 304 -47 305 -27
<< ndcontact >>
rect -204 -5 -200 5
rect -196 -5 -192 5
rect -168 -5 -164 5
rect -160 -5 -156 5
rect -152 -5 -148 5
rect -124 -5 -120 5
rect -116 -5 -112 5
rect -108 -5 -104 5
rect -73 -5 -69 5
rect -65 -5 -61 5
rect 9 -5 13 5
rect 17 -5 21 5
rect 45 -5 49 5
rect 53 -5 57 5
rect 61 -5 65 5
rect 89 -5 93 5
rect 97 -5 101 5
rect 105 -5 109 5
rect 140 -5 144 5
rect 148 -5 152 5
rect 297 -7 301 13
rect 305 -7 309 13
rect 506 -12 510 0
rect 524 -12 528 0
rect 546 -1 550 5
rect 554 -1 558 5
rect 260 -59 264 -39
rect 268 -59 272 -39
rect 330 -54 334 -34
rect 338 -54 342 -34
rect 373 -60 377 -40
rect 381 -60 385 -40
<< pdcontact >>
rect -200 27 -196 52
rect -192 27 -188 52
rect -184 27 -180 52
rect -162 27 -158 52
rect -154 27 -150 52
rect -118 27 -114 52
rect -110 27 -106 52
rect -73 27 -69 52
rect -65 27 -61 52
rect 13 27 17 52
rect 21 27 25 52
rect 29 27 33 52
rect 51 27 55 52
rect 59 27 63 52
rect 95 27 99 52
rect 103 27 107 52
rect 140 27 144 52
rect 148 27 152 52
rect 260 -19 264 21
rect 268 -19 272 21
rect 506 20 510 32
rect 515 20 519 32
rect 524 20 528 32
rect 330 -14 334 6
rect 338 -14 342 6
rect 373 -20 377 20
rect 381 -20 385 20
rect 546 19 550 31
rect 554 19 558 31
rect 297 -47 301 -27
rect 305 -47 309 -27
<< polysilicon >>
rect -195 52 -193 55
rect -187 52 -185 55
rect -157 52 -155 55
rect -113 52 -111 55
rect -68 52 -66 55
rect 18 52 20 55
rect 26 52 28 55
rect 56 52 58 55
rect 100 52 102 55
rect 145 52 147 55
rect 511 32 513 35
rect 521 32 523 35
rect -195 20 -193 27
rect -200 16 -193 20
rect -199 5 -197 16
rect -187 8 -185 27
rect -157 19 -155 27
rect -113 19 -111 27
rect -163 17 -155 19
rect -119 17 -111 19
rect -163 5 -161 17
rect -155 5 -153 14
rect -119 5 -117 17
rect -111 5 -109 14
rect -68 5 -66 27
rect 18 20 20 27
rect 13 16 20 20
rect 14 5 16 16
rect 26 8 28 27
rect 56 19 58 27
rect 100 19 102 27
rect 50 17 58 19
rect 94 17 102 19
rect 50 5 52 17
rect 58 5 60 14
rect 94 5 96 17
rect 102 5 104 14
rect 145 5 147 27
rect 265 21 267 25
rect -199 -8 -197 -5
rect -163 -8 -161 -5
rect -155 -8 -153 -5
rect -119 -8 -117 -5
rect -111 -8 -109 -5
rect -68 -8 -66 -5
rect 14 -8 16 -5
rect 50 -8 52 -5
rect 58 -8 60 -5
rect 94 -8 96 -5
rect 102 -8 104 -5
rect 145 -8 147 -5
rect 378 20 380 24
rect 551 31 553 34
rect 302 13 304 20
rect 335 6 337 20
rect 302 -10 304 -7
rect 335 -17 337 -14
rect 265 -39 267 -19
rect 511 0 513 20
rect 521 0 523 20
rect 551 5 553 19
rect 551 -4 553 -1
rect 511 -15 513 -12
rect 521 -15 523 -12
rect 302 -27 304 -24
rect 335 -34 337 -31
rect 265 -62 267 -59
rect 302 -61 304 -47
rect 378 -40 380 -20
rect 335 -61 337 -54
rect 378 -63 380 -60
<< polycontact >>
rect -204 16 -200 20
rect -191 8 -187 12
rect -168 8 -163 13
rect -153 8 -148 12
rect -124 8 -119 13
rect -72 13 -68 18
rect -109 8 -104 12
rect 9 16 13 20
rect 22 8 26 12
rect 45 8 50 13
rect 60 8 65 12
rect 89 8 94 13
rect 141 13 145 18
rect 104 8 109 12
rect 301 20 305 25
rect 334 20 338 25
rect 261 -36 265 -31
rect 507 9 511 13
rect 517 3 521 7
rect 547 8 551 12
rect 374 -37 378 -32
rect 301 -66 305 -61
rect 334 -66 338 -61
<< metal1 >>
rect -206 58 498 62
rect -200 52 -196 58
rect -162 52 -158 58
rect -118 52 -114 58
rect -73 52 -69 58
rect 13 52 17 58
rect 51 52 55 58
rect 95 52 99 58
rect 140 52 144 58
rect 232 57 498 58
rect -150 27 -137 52
rect -106 27 -93 52
rect 63 27 76 52
rect 107 27 120 52
rect -211 16 -204 20
rect -184 19 -180 27
rect -184 16 -144 19
rect -194 8 -191 12
rect -184 5 -180 16
rect -172 8 -168 13
rect -148 8 -144 16
rect -140 13 -137 27
rect -96 18 -93 27
rect -96 13 -72 18
rect -65 17 -61 27
rect -140 8 -124 13
rect -104 8 -100 12
rect -140 5 -137 8
rect -96 5 -93 13
rect -65 12 -52 17
rect -65 5 -61 12
rect 2 16 9 20
rect 29 19 33 27
rect 29 16 69 19
rect 19 8 22 12
rect 29 5 33 16
rect 41 8 45 13
rect 65 8 69 16
rect 73 13 76 27
rect 117 18 120 27
rect 117 13 141 18
rect 148 17 152 27
rect 260 21 264 57
rect 73 8 89 13
rect 109 8 113 12
rect 73 5 76 8
rect 117 5 120 13
rect 148 12 161 17
rect 148 5 152 12
rect -192 -5 -180 5
rect -148 -5 -137 5
rect -104 -5 -93 5
rect 21 -5 33 5
rect 65 -5 76 5
rect 109 -5 120 5
rect -204 -10 -200 -5
rect -168 -10 -164 -5
rect -124 -10 -120 -5
rect -73 -10 -69 -5
rect 9 -10 13 -5
rect 45 -10 49 -5
rect 89 -10 93 -5
rect 140 -10 144 -5
rect -205 -14 152 -10
rect 148 -99 152 -14
rect 285 -11 290 44
rect 301 25 305 32
rect 334 25 338 32
rect 373 20 377 57
rect 460 37 466 44
rect 493 41 498 57
rect 493 40 543 41
rect 493 38 564 40
rect 393 32 474 37
rect 297 -11 301 -7
rect 285 -15 301 -11
rect 251 -36 261 -31
rect 268 -32 272 -19
rect 297 -27 301 -15
rect 268 -37 281 -32
rect 268 -39 272 -37
rect 305 -12 309 -7
rect 305 -16 322 -12
rect 305 -27 309 -16
rect 318 -26 322 -16
rect 330 -26 334 -14
rect 318 -31 334 -26
rect 260 -98 264 -59
rect 301 -79 305 -66
rect 318 -92 324 -31
rect 330 -34 334 -31
rect 338 -27 342 -14
rect 338 -31 359 -27
rect 338 -34 342 -31
rect 353 -32 359 -31
rect 353 -37 363 -32
rect 369 -37 374 -32
rect 381 -33 385 -20
rect 423 6 432 19
rect 471 12 474 32
rect 506 32 509 38
rect 525 32 528 38
rect 540 37 564 38
rect 546 31 549 37
rect 515 17 518 20
rect 515 14 528 17
rect 471 9 507 12
rect 525 11 528 14
rect 525 8 547 11
rect 555 11 558 19
rect 555 8 567 11
rect 423 3 517 6
rect 381 -38 398 -33
rect 381 -40 385 -38
rect 334 -79 338 -66
rect 373 -98 377 -60
rect 423 -78 431 3
rect 525 0 528 8
rect 555 5 558 8
rect 546 -5 549 -1
rect 536 -8 564 -5
rect 506 -18 509 -12
rect 536 -18 540 -8
rect 441 -21 540 -18
rect 441 -98 452 -21
rect 232 -99 452 -98
rect 148 -106 452 -99
<< m2contact >>
rect -52 11 -41 18
rect 285 44 291 49
rect 161 11 172 18
rect 301 32 306 37
rect 333 32 338 37
rect 457 44 467 51
rect 385 32 393 37
rect 246 -36 251 -31
rect 281 -37 287 -32
rect 301 -84 306 -79
rect 422 19 433 25
rect 363 -37 369 -32
rect 398 -38 404 -33
rect 334 -84 339 -79
rect 423 -84 431 -78
<< metal2 >>
rect 187 80 191 81
rect 187 76 465 80
rect -26 65 169 69
rect -26 17 -22 65
rect -41 12 -22 17
rect 187 17 191 76
rect 230 67 430 71
rect 291 44 404 49
rect 172 12 191 17
rect 246 32 301 37
rect 306 32 333 37
rect 338 32 385 37
rect 246 -31 250 32
rect 281 -79 287 -37
rect 363 -78 369 -37
rect 398 -33 404 44
rect 424 25 430 67
rect 460 51 465 76
rect 280 -84 301 -79
rect 306 -84 334 -79
rect 339 -84 353 -79
rect 363 -84 423 -78
<< m3contact >>
rect 169 64 182 70
rect 220 65 230 71
<< metal3 >>
rect 182 65 220 70
<< labels >>
rlabel metal1 562 8 567 11 1 g0
rlabel metal1 500 3 503 6 1 b0_reg
rlabel metal1 500 9 504 12 1 a0_reg
rlabel metal1 560 -7 560 -7 1 gnd!
rlabel metal1 554 38 554 38 5 vdd!
rlabel metal1 534 8 534 11 7 out
rlabel metal1 524 -20 524 -20 1 gnd!
rlabel metal1 524 40 524 40 5 vdd!
rlabel metal1 457 32 472 37 1 a0_reg
rlabel metal1 423 -19 431 -3 1 b0_reg
rlabel metal1 318 -91 324 -85 1 p0
rlabel metal1 341 57 455 62 1 vdd
rlabel metal1 317 -105 431 -99 1 gnd
rlabel metal1 19 9 21 11 1 clk
rlabel metal1 17 -12 20 -11 1 gnd
rlabel metal1 23 60 25 61 5 vdd
rlabel metal1 42 9 43 11 1 clk
rlabel metal1 110 9 112 11 1 clk
rlabel metal1 154 14 157 16 1 a0_reg
rlabel metal1 4 17 6 19 3 a0
rlabel metal1 -103 9 -101 11 1 clk
rlabel metal1 -171 9 -170 11 1 clk
rlabel metal1 -190 60 -188 61 5 vdd
rlabel metal1 -196 -12 -193 -11 1 gnd
rlabel metal1 -194 9 -192 11 1 clk
rlabel metal1 -209 17 -207 19 3 b0
rlabel metal1 -59 14 -56 16 1 b0_reg
<< end >>
