.include TSMC_180nm.txt
.param SUPPLY=1.8

.global gnd vdd
.option scale=0.09u
Vdd    vdd gnd 'SUPPLY'
vin    in 0 pulse 0 1.8 0ns 0ns 0ns 10ns 20ns

M1000 op in vdd w_0_6# CMOSP w=12 l=2
+  ad=60 pd=34 as=60 ps=34
M1001 op in gnd Gnd CMOSN w=6 l=2
+  ad=30 pd=22 as=30 ps=22
C0 vdd w_0_6# 0.06fF
C1 gnd op 0.10fF
C2 op in 0.04fF
C3 gnd in 0.05fF
C4 vdd op 0.15fF
C5 vdd in 0.02fF
C6 w_0_6# op 0.03fF
C7 w_0_6# in 0.06fF
C8 gnd Gnd 0.09fF
C9 op Gnd 0.05fF
C10 vdd Gnd 0.03fF
C11 in Gnd 0.14fF
C12 w_0_6# Gnd 0.58fF


    .tran 0.1n 200n
    .control
    run
     set curplottitle  = "Eswar-2023102011"
    plot 5+v(in)  v(op)
    .endc
