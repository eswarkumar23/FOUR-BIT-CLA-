magic
tech scmos
timestamp 1732886045
<< nwell >>
rect -1520 294 -1488 331
rect -1482 294 -1456 331
rect -1438 294 -1412 331
rect -1393 294 -1367 331
rect -1307 294 -1275 331
rect -1269 294 -1243 331
rect -1225 294 -1199 331
rect -1180 294 -1154 331
rect -1060 244 -1035 301
rect -1023 216 -998 256
rect -990 249 -965 289
rect -947 243 -922 300
rect -814 287 -780 311
rect -774 286 -750 310
rect -631 256 -599 293
rect -593 256 -567 293
rect -549 256 -523 293
rect -504 256 -478 293
rect -379 144 -355 206
rect -290 144 -266 206
rect -227 144 -203 206
rect -172 144 -148 206
rect -121 181 -97 233
rect -83 181 -59 233
rect -39 181 -15 233
rect -1 181 23 233
rect 248 111 273 168
rect 285 83 310 123
rect 318 116 343 156
rect 361 110 386 167
rect 590 143 622 180
rect 628 143 654 180
rect 672 143 698 180
rect 717 143 743 180
rect -1505 -35 -1473 2
rect -1467 -35 -1441 2
rect -1423 -35 -1397 2
rect -1378 -35 -1352 2
rect -1292 -35 -1260 2
rect -1254 -35 -1228 2
rect -1210 -35 -1184 2
rect -1165 -35 -1139 2
rect -1045 -85 -1020 -28
rect -1008 -113 -983 -73
rect -975 -80 -950 -40
rect -932 -86 -907 -29
rect -799 -42 -765 -18
rect -759 -43 -735 -19
rect -597 -36 -573 -12
rect 238 -197 263 -140
rect 275 -225 300 -185
rect 308 -192 333 -152
rect 351 -198 376 -141
rect 580 -165 612 -128
rect 618 -165 644 -128
rect 662 -165 688 -128
rect 707 -165 733 -128
rect -1481 -302 -1449 -265
rect -1443 -302 -1417 -265
rect -1399 -302 -1373 -265
rect -1354 -302 -1328 -265
rect -1268 -302 -1236 -265
rect -1230 -302 -1204 -265
rect -1186 -302 -1160 -265
rect -1141 -302 -1115 -265
rect -1021 -352 -996 -295
rect -984 -380 -959 -340
rect -951 -347 -926 -307
rect -908 -353 -883 -296
rect -775 -309 -741 -285
rect -735 -310 -711 -286
rect 262 -456 287 -399
rect 299 -484 324 -444
rect 332 -451 357 -411
rect 375 -457 400 -400
rect 604 -424 636 -387
rect 642 -424 668 -387
rect 686 -424 712 -387
rect 731 -424 757 -387
rect -1452 -612 -1420 -575
rect -1414 -612 -1388 -575
rect -1370 -612 -1344 -575
rect -1325 -612 -1299 -575
rect -1239 -612 -1207 -575
rect -1201 -612 -1175 -575
rect -1157 -612 -1131 -575
rect -1112 -612 -1086 -575
rect -992 -662 -967 -605
rect -955 -690 -930 -650
rect -922 -657 -897 -617
rect -879 -663 -854 -606
rect -746 -619 -712 -595
rect -706 -620 -682 -596
rect 283 -762 308 -705
rect 320 -790 345 -750
rect 353 -757 378 -717
rect 396 -763 421 -706
rect 625 -730 657 -693
rect 663 -730 689 -693
rect 707 -730 733 -693
rect 752 -730 778 -693
rect 690 -970 722 -933
rect 728 -970 754 -933
rect 772 -970 798 -933
rect 817 -970 843 -933
<< ntransistor >>
rect -1513 268 -1511 278
rect -1477 268 -1475 278
rect -1469 268 -1467 278
rect -1433 268 -1431 278
rect -1425 268 -1423 278
rect -1382 268 -1380 278
rect -1300 268 -1298 278
rect -1264 268 -1262 278
rect -1256 268 -1254 278
rect -1220 268 -1218 278
rect -1212 268 -1210 278
rect -1169 268 -1167 278
rect -1012 266 -1010 286
rect -803 261 -801 273
rect -793 261 -791 273
rect -763 272 -761 278
rect -1049 214 -1047 234
rect -979 219 -977 239
rect -936 213 -934 233
rect -624 230 -622 240
rect -588 230 -586 240
rect -580 230 -578 240
rect -544 230 -542 240
rect -536 230 -534 240
rect -493 230 -491 240
rect -110 149 -108 169
rect -72 149 -70 169
rect -28 149 -26 169
rect 10 149 12 169
rect 296 133 298 153
rect -153 11 -151 111
rect -75 10 -73 110
rect 259 81 261 101
rect 329 86 331 106
rect 597 117 599 127
rect 633 117 635 127
rect 641 117 643 127
rect 677 117 679 127
rect 685 117 687 127
rect 728 117 730 127
rect 372 80 374 100
rect -1498 -61 -1496 -51
rect -1462 -61 -1460 -51
rect -1454 -61 -1452 -51
rect -1418 -61 -1416 -51
rect -1410 -61 -1408 -51
rect -1367 -61 -1365 -51
rect -1285 -61 -1283 -51
rect -1249 -61 -1247 -51
rect -1241 -61 -1239 -51
rect -1205 -61 -1203 -51
rect -1197 -61 -1195 -51
rect -1154 -61 -1152 -51
rect -997 -63 -995 -43
rect -586 -50 -584 -44
rect -788 -68 -786 -56
rect -778 -68 -776 -56
rect -748 -57 -746 -51
rect -1034 -115 -1032 -95
rect -964 -110 -962 -90
rect -921 -116 -919 -96
rect -208 -127 -206 -27
rect -145 -128 -143 -28
rect -271 -272 -269 -172
rect -200 -272 -198 -172
rect 286 -175 288 -155
rect 249 -227 251 -207
rect 319 -222 321 -202
rect 587 -191 589 -181
rect 623 -191 625 -181
rect 631 -191 633 -181
rect 667 -191 669 -181
rect 675 -191 677 -181
rect 718 -191 720 -181
rect 362 -228 364 -208
rect -1474 -328 -1472 -318
rect -1438 -328 -1436 -318
rect -1430 -328 -1428 -318
rect -1394 -328 -1392 -318
rect -1386 -328 -1384 -318
rect -1343 -328 -1341 -318
rect -1261 -328 -1259 -318
rect -1225 -328 -1223 -318
rect -1217 -328 -1215 -318
rect -1181 -328 -1179 -318
rect -1173 -328 -1171 -318
rect -1130 -328 -1128 -318
rect -973 -330 -971 -310
rect -764 -335 -762 -323
rect -754 -335 -752 -323
rect -724 -324 -722 -318
rect -1010 -382 -1008 -362
rect -940 -377 -938 -357
rect -897 -383 -895 -363
rect -360 -420 -358 -320
rect -263 -420 -261 -320
rect 310 -434 312 -414
rect -352 -565 -350 -465
rect 273 -486 275 -466
rect 343 -481 345 -461
rect 611 -450 613 -440
rect 647 -450 649 -440
rect 655 -450 657 -440
rect 691 -450 693 -440
rect 699 -450 701 -440
rect 742 -450 744 -440
rect 386 -487 388 -467
rect -1445 -638 -1443 -628
rect -1409 -638 -1407 -628
rect -1401 -638 -1399 -628
rect -1365 -638 -1363 -628
rect -1357 -638 -1355 -628
rect -1314 -638 -1312 -628
rect -1232 -638 -1230 -628
rect -1196 -638 -1194 -628
rect -1188 -638 -1186 -628
rect -1152 -638 -1150 -628
rect -1144 -638 -1142 -628
rect -1101 -638 -1099 -628
rect -944 -640 -942 -620
rect -735 -645 -733 -633
rect -725 -645 -723 -633
rect -695 -634 -693 -628
rect -981 -692 -979 -672
rect -911 -687 -909 -667
rect -868 -693 -866 -673
rect -344 -698 -342 -598
rect 331 -740 333 -720
rect 294 -792 296 -772
rect 364 -787 366 -767
rect 632 -756 634 -746
rect 668 -756 670 -746
rect 676 -756 678 -746
rect 712 -756 714 -746
rect 720 -756 722 -746
rect 763 -756 765 -746
rect 407 -793 409 -773
rect 697 -996 699 -986
rect 733 -996 735 -986
rect 741 -996 743 -986
rect 777 -996 779 -986
rect 785 -996 787 -986
rect 828 -996 830 -986
<< ptransistor >>
rect -1509 300 -1507 325
rect -1501 300 -1499 325
rect -1471 300 -1469 325
rect -1427 300 -1425 325
rect -1382 300 -1380 325
rect -1296 300 -1294 325
rect -1288 300 -1286 325
rect -1258 300 -1256 325
rect -1214 300 -1212 325
rect -1169 300 -1167 325
rect -1049 254 -1047 294
rect -803 293 -801 305
rect -793 293 -791 305
rect -979 259 -977 279
rect -936 253 -934 293
rect -763 292 -761 304
rect -620 262 -618 287
rect -612 262 -610 287
rect -582 262 -580 287
rect -538 262 -536 287
rect -493 262 -491 287
rect -1012 226 -1010 246
rect -368 150 -366 200
rect -279 150 -277 200
rect -216 150 -214 200
rect -161 150 -159 200
rect -110 187 -108 227
rect -72 187 -70 227
rect -28 187 -26 227
rect 10 187 12 227
rect 259 121 261 161
rect 329 126 331 146
rect 372 120 374 160
rect 601 149 603 174
rect 609 149 611 174
rect 639 149 641 174
rect 683 149 685 174
rect 728 149 730 174
rect 296 93 298 113
rect -1494 -29 -1492 -4
rect -1486 -29 -1484 -4
rect -1456 -29 -1454 -4
rect -1412 -29 -1410 -4
rect -1367 -29 -1365 -4
rect -1281 -29 -1279 -4
rect -1273 -29 -1271 -4
rect -1243 -29 -1241 -4
rect -1199 -29 -1197 -4
rect -1154 -29 -1152 -4
rect -1034 -75 -1032 -35
rect -788 -36 -786 -24
rect -778 -36 -776 -24
rect -964 -70 -962 -50
rect -921 -76 -919 -36
rect -748 -37 -746 -25
rect -586 -30 -584 -18
rect -997 -103 -995 -83
rect -1470 -296 -1468 -271
rect -1462 -296 -1460 -271
rect -1432 -296 -1430 -271
rect -1388 -296 -1386 -271
rect -1343 -296 -1341 -271
rect -1257 -296 -1255 -271
rect -1249 -296 -1247 -271
rect -1219 -296 -1217 -271
rect -1175 -296 -1173 -271
rect -1130 -296 -1128 -271
rect 249 -187 251 -147
rect 319 -182 321 -162
rect 362 -188 364 -148
rect 591 -159 593 -134
rect 599 -159 601 -134
rect 629 -159 631 -134
rect 673 -159 675 -134
rect 718 -159 720 -134
rect 286 -215 288 -195
rect -1010 -342 -1008 -302
rect -764 -303 -762 -291
rect -754 -303 -752 -291
rect -940 -337 -938 -317
rect -897 -343 -895 -303
rect -724 -304 -722 -292
rect -973 -370 -971 -350
rect 273 -446 275 -406
rect 343 -441 345 -421
rect 386 -447 388 -407
rect 615 -418 617 -393
rect 623 -418 625 -393
rect 653 -418 655 -393
rect 697 -418 699 -393
rect 742 -418 744 -393
rect 310 -474 312 -454
rect -1441 -606 -1439 -581
rect -1433 -606 -1431 -581
rect -1403 -606 -1401 -581
rect -1359 -606 -1357 -581
rect -1314 -606 -1312 -581
rect -1228 -606 -1226 -581
rect -1220 -606 -1218 -581
rect -1190 -606 -1188 -581
rect -1146 -606 -1144 -581
rect -1101 -606 -1099 -581
rect -981 -652 -979 -612
rect -735 -613 -733 -601
rect -725 -613 -723 -601
rect -911 -647 -909 -627
rect -868 -653 -866 -613
rect -695 -614 -693 -602
rect -944 -680 -942 -660
rect 294 -752 296 -712
rect 364 -747 366 -727
rect 407 -753 409 -713
rect 636 -724 638 -699
rect 644 -724 646 -699
rect 674 -724 676 -699
rect 718 -724 720 -699
rect 763 -724 765 -699
rect 331 -780 333 -760
rect 701 -964 703 -939
rect 709 -964 711 -939
rect 739 -964 741 -939
rect 783 -964 785 -939
rect 828 -964 830 -939
<< ndiffusion >>
rect -1514 268 -1513 278
rect -1511 268 -1510 278
rect -1478 268 -1477 278
rect -1475 268 -1474 278
rect -1470 268 -1469 278
rect -1467 268 -1466 278
rect -1434 268 -1433 278
rect -1431 268 -1430 278
rect -1426 268 -1425 278
rect -1423 268 -1422 278
rect -1383 268 -1382 278
rect -1380 268 -1379 278
rect -1301 268 -1300 278
rect -1298 268 -1297 278
rect -1265 268 -1264 278
rect -1262 268 -1261 278
rect -1257 268 -1256 278
rect -1254 268 -1253 278
rect -1221 268 -1220 278
rect -1218 268 -1217 278
rect -1213 268 -1212 278
rect -1210 268 -1209 278
rect -1170 268 -1169 278
rect -1167 268 -1166 278
rect -1013 266 -1012 286
rect -1010 266 -1009 286
rect -804 261 -803 273
rect -801 261 -793 273
rect -791 261 -790 273
rect -764 272 -763 278
rect -761 272 -760 278
rect -1050 214 -1049 234
rect -1047 214 -1046 234
rect -980 219 -979 239
rect -977 219 -976 239
rect -937 213 -936 233
rect -934 213 -933 233
rect -625 230 -624 240
rect -622 230 -621 240
rect -589 230 -588 240
rect -586 230 -585 240
rect -581 230 -580 240
rect -578 230 -577 240
rect -545 230 -544 240
rect -542 230 -541 240
rect -537 230 -536 240
rect -534 230 -533 240
rect -494 230 -493 240
rect -491 230 -490 240
rect -111 149 -110 169
rect -108 149 -107 169
rect -73 149 -72 169
rect -70 149 -69 169
rect -29 149 -28 169
rect -26 149 -25 169
rect 9 149 10 169
rect 12 149 13 169
rect 295 133 296 153
rect 298 133 299 153
rect -154 11 -153 111
rect -151 11 -150 111
rect -76 10 -75 110
rect -73 10 -72 110
rect 258 81 259 101
rect 261 81 262 101
rect 328 86 329 106
rect 331 86 332 106
rect 596 117 597 127
rect 599 117 600 127
rect 632 117 633 127
rect 635 117 636 127
rect 640 117 641 127
rect 643 117 644 127
rect 676 117 677 127
rect 679 117 680 127
rect 684 117 685 127
rect 687 117 688 127
rect 727 117 728 127
rect 730 117 731 127
rect 371 80 372 100
rect 374 80 375 100
rect -1499 -61 -1498 -51
rect -1496 -61 -1495 -51
rect -1463 -61 -1462 -51
rect -1460 -61 -1459 -51
rect -1455 -61 -1454 -51
rect -1452 -61 -1451 -51
rect -1419 -61 -1418 -51
rect -1416 -61 -1415 -51
rect -1411 -61 -1410 -51
rect -1408 -61 -1407 -51
rect -1368 -61 -1367 -51
rect -1365 -61 -1364 -51
rect -1286 -61 -1285 -51
rect -1283 -61 -1282 -51
rect -1250 -61 -1249 -51
rect -1247 -61 -1246 -51
rect -1242 -61 -1241 -51
rect -1239 -61 -1238 -51
rect -1206 -61 -1205 -51
rect -1203 -61 -1202 -51
rect -1198 -61 -1197 -51
rect -1195 -61 -1194 -51
rect -1155 -61 -1154 -51
rect -1152 -61 -1151 -51
rect -998 -63 -997 -43
rect -995 -63 -994 -43
rect -587 -50 -586 -44
rect -584 -50 -583 -44
rect -789 -68 -788 -56
rect -786 -68 -778 -56
rect -776 -68 -775 -56
rect -749 -57 -748 -51
rect -746 -57 -745 -51
rect -1035 -115 -1034 -95
rect -1032 -115 -1031 -95
rect -965 -110 -964 -90
rect -962 -110 -961 -90
rect -922 -116 -921 -96
rect -919 -116 -918 -96
rect -209 -127 -208 -27
rect -206 -127 -205 -27
rect -146 -128 -145 -28
rect -143 -128 -142 -28
rect -272 -272 -271 -172
rect -269 -272 -268 -172
rect -201 -272 -200 -172
rect -198 -272 -197 -172
rect 285 -175 286 -155
rect 288 -175 289 -155
rect 248 -227 249 -207
rect 251 -227 252 -207
rect 318 -222 319 -202
rect 321 -222 322 -202
rect 586 -191 587 -181
rect 589 -191 590 -181
rect 622 -191 623 -181
rect 625 -191 626 -181
rect 630 -191 631 -181
rect 633 -191 634 -181
rect 666 -191 667 -181
rect 669 -191 670 -181
rect 674 -191 675 -181
rect 677 -191 678 -181
rect 717 -191 718 -181
rect 720 -191 721 -181
rect 361 -228 362 -208
rect 364 -228 365 -208
rect -1475 -328 -1474 -318
rect -1472 -328 -1471 -318
rect -1439 -328 -1438 -318
rect -1436 -328 -1435 -318
rect -1431 -328 -1430 -318
rect -1428 -328 -1427 -318
rect -1395 -328 -1394 -318
rect -1392 -328 -1391 -318
rect -1387 -328 -1386 -318
rect -1384 -328 -1383 -318
rect -1344 -328 -1343 -318
rect -1341 -328 -1340 -318
rect -1262 -328 -1261 -318
rect -1259 -328 -1258 -318
rect -1226 -328 -1225 -318
rect -1223 -328 -1222 -318
rect -1218 -328 -1217 -318
rect -1215 -328 -1214 -318
rect -1182 -328 -1181 -318
rect -1179 -328 -1178 -318
rect -1174 -328 -1173 -318
rect -1171 -328 -1170 -318
rect -1131 -328 -1130 -318
rect -1128 -328 -1127 -318
rect -974 -330 -973 -310
rect -971 -330 -970 -310
rect -765 -335 -764 -323
rect -762 -335 -754 -323
rect -752 -335 -751 -323
rect -725 -324 -724 -318
rect -722 -324 -721 -318
rect -1011 -382 -1010 -362
rect -1008 -382 -1007 -362
rect -941 -377 -940 -357
rect -938 -377 -937 -357
rect -898 -383 -897 -363
rect -895 -383 -894 -363
rect -361 -420 -360 -320
rect -358 -420 -357 -320
rect -264 -420 -263 -320
rect -261 -420 -260 -320
rect 309 -434 310 -414
rect 312 -434 313 -414
rect -353 -565 -352 -465
rect -350 -565 -349 -465
rect 272 -486 273 -466
rect 275 -486 276 -466
rect 342 -481 343 -461
rect 345 -481 346 -461
rect 610 -450 611 -440
rect 613 -450 614 -440
rect 646 -450 647 -440
rect 649 -450 650 -440
rect 654 -450 655 -440
rect 657 -450 658 -440
rect 690 -450 691 -440
rect 693 -450 694 -440
rect 698 -450 699 -440
rect 701 -450 702 -440
rect 741 -450 742 -440
rect 744 -450 745 -440
rect 385 -487 386 -467
rect 388 -487 389 -467
rect -1446 -638 -1445 -628
rect -1443 -638 -1442 -628
rect -1410 -638 -1409 -628
rect -1407 -638 -1406 -628
rect -1402 -638 -1401 -628
rect -1399 -638 -1398 -628
rect -1366 -638 -1365 -628
rect -1363 -638 -1362 -628
rect -1358 -638 -1357 -628
rect -1355 -638 -1354 -628
rect -1315 -638 -1314 -628
rect -1312 -638 -1311 -628
rect -1233 -638 -1232 -628
rect -1230 -638 -1229 -628
rect -1197 -638 -1196 -628
rect -1194 -638 -1193 -628
rect -1189 -638 -1188 -628
rect -1186 -638 -1185 -628
rect -1153 -638 -1152 -628
rect -1150 -638 -1149 -628
rect -1145 -638 -1144 -628
rect -1142 -638 -1141 -628
rect -1102 -638 -1101 -628
rect -1099 -638 -1098 -628
rect -945 -640 -944 -620
rect -942 -640 -941 -620
rect -736 -645 -735 -633
rect -733 -645 -725 -633
rect -723 -645 -722 -633
rect -696 -634 -695 -628
rect -693 -634 -692 -628
rect -982 -692 -981 -672
rect -979 -692 -978 -672
rect -912 -687 -911 -667
rect -909 -687 -908 -667
rect -869 -693 -868 -673
rect -866 -693 -865 -673
rect -345 -698 -344 -598
rect -342 -698 -341 -598
rect 330 -740 331 -720
rect 333 -740 334 -720
rect 293 -792 294 -772
rect 296 -792 297 -772
rect 363 -787 364 -767
rect 366 -787 367 -767
rect 631 -756 632 -746
rect 634 -756 635 -746
rect 667 -756 668 -746
rect 670 -756 671 -746
rect 675 -756 676 -746
rect 678 -756 679 -746
rect 711 -756 712 -746
rect 714 -756 715 -746
rect 719 -756 720 -746
rect 722 -756 723 -746
rect 762 -756 763 -746
rect 765 -756 766 -746
rect 406 -793 407 -773
rect 409 -793 410 -773
rect 696 -996 697 -986
rect 699 -996 700 -986
rect 732 -996 733 -986
rect 735 -996 736 -986
rect 740 -996 741 -986
rect 743 -996 744 -986
rect 776 -996 777 -986
rect 779 -996 780 -986
rect 784 -996 785 -986
rect 787 -996 788 -986
rect 827 -996 828 -986
rect 830 -996 831 -986
<< pdiffusion >>
rect -1510 300 -1509 325
rect -1507 300 -1506 325
rect -1502 300 -1501 325
rect -1499 300 -1498 325
rect -1472 300 -1471 325
rect -1469 300 -1468 325
rect -1428 300 -1427 325
rect -1425 300 -1424 325
rect -1383 300 -1382 325
rect -1380 300 -1379 325
rect -1297 300 -1296 325
rect -1294 300 -1293 325
rect -1289 300 -1288 325
rect -1286 300 -1285 325
rect -1259 300 -1258 325
rect -1256 300 -1255 325
rect -1215 300 -1214 325
rect -1212 300 -1211 325
rect -1170 300 -1169 325
rect -1167 300 -1166 325
rect -1050 254 -1049 294
rect -1047 254 -1046 294
rect -804 293 -803 305
rect -801 293 -799 305
rect -795 293 -793 305
rect -791 293 -790 305
rect -980 259 -979 279
rect -977 259 -976 279
rect -937 253 -936 293
rect -934 253 -933 293
rect -764 292 -763 304
rect -761 292 -760 304
rect -621 262 -620 287
rect -618 262 -617 287
rect -613 262 -612 287
rect -610 262 -609 287
rect -583 262 -582 287
rect -580 262 -579 287
rect -539 262 -538 287
rect -536 262 -535 287
rect -494 262 -493 287
rect -491 262 -490 287
rect -1013 226 -1012 246
rect -1010 226 -1009 246
rect -369 150 -368 200
rect -366 150 -365 200
rect -280 150 -279 200
rect -277 150 -276 200
rect -217 150 -216 200
rect -214 150 -213 200
rect -162 150 -161 200
rect -159 150 -158 200
rect -111 187 -110 227
rect -108 187 -107 227
rect -73 187 -72 227
rect -70 187 -69 227
rect -29 187 -28 227
rect -26 187 -25 227
rect 9 187 10 227
rect 12 187 13 227
rect 258 121 259 161
rect 261 121 262 161
rect 328 126 329 146
rect 331 126 332 146
rect 371 120 372 160
rect 374 120 375 160
rect 600 149 601 174
rect 603 149 604 174
rect 608 149 609 174
rect 611 149 612 174
rect 638 149 639 174
rect 641 149 642 174
rect 682 149 683 174
rect 685 149 686 174
rect 727 149 728 174
rect 730 149 731 174
rect 295 93 296 113
rect 298 93 299 113
rect -1495 -29 -1494 -4
rect -1492 -29 -1491 -4
rect -1487 -29 -1486 -4
rect -1484 -29 -1483 -4
rect -1457 -29 -1456 -4
rect -1454 -29 -1453 -4
rect -1413 -29 -1412 -4
rect -1410 -29 -1409 -4
rect -1368 -29 -1367 -4
rect -1365 -29 -1364 -4
rect -1282 -29 -1281 -4
rect -1279 -29 -1278 -4
rect -1274 -29 -1273 -4
rect -1271 -29 -1270 -4
rect -1244 -29 -1243 -4
rect -1241 -29 -1240 -4
rect -1200 -29 -1199 -4
rect -1197 -29 -1196 -4
rect -1155 -29 -1154 -4
rect -1152 -29 -1151 -4
rect -1035 -75 -1034 -35
rect -1032 -75 -1031 -35
rect -789 -36 -788 -24
rect -786 -36 -784 -24
rect -780 -36 -778 -24
rect -776 -36 -775 -24
rect -965 -70 -964 -50
rect -962 -70 -961 -50
rect -922 -76 -921 -36
rect -919 -76 -918 -36
rect -749 -37 -748 -25
rect -746 -37 -745 -25
rect -587 -30 -586 -18
rect -584 -30 -583 -18
rect -998 -103 -997 -83
rect -995 -103 -994 -83
rect -1471 -296 -1470 -271
rect -1468 -296 -1467 -271
rect -1463 -296 -1462 -271
rect -1460 -296 -1459 -271
rect -1433 -296 -1432 -271
rect -1430 -296 -1429 -271
rect -1389 -296 -1388 -271
rect -1386 -296 -1385 -271
rect -1344 -296 -1343 -271
rect -1341 -296 -1340 -271
rect -1258 -296 -1257 -271
rect -1255 -296 -1254 -271
rect -1250 -296 -1249 -271
rect -1247 -296 -1246 -271
rect -1220 -296 -1219 -271
rect -1217 -296 -1216 -271
rect -1176 -296 -1175 -271
rect -1173 -296 -1172 -271
rect -1131 -296 -1130 -271
rect -1128 -296 -1127 -271
rect 248 -187 249 -147
rect 251 -187 252 -147
rect 318 -182 319 -162
rect 321 -182 322 -162
rect 361 -188 362 -148
rect 364 -188 365 -148
rect 590 -159 591 -134
rect 593 -159 594 -134
rect 598 -159 599 -134
rect 601 -159 602 -134
rect 628 -159 629 -134
rect 631 -159 632 -134
rect 672 -159 673 -134
rect 675 -159 676 -134
rect 717 -159 718 -134
rect 720 -159 721 -134
rect 285 -215 286 -195
rect 288 -215 289 -195
rect -1011 -342 -1010 -302
rect -1008 -342 -1007 -302
rect -765 -303 -764 -291
rect -762 -303 -760 -291
rect -756 -303 -754 -291
rect -752 -303 -751 -291
rect -941 -337 -940 -317
rect -938 -337 -937 -317
rect -898 -343 -897 -303
rect -895 -343 -894 -303
rect -725 -304 -724 -292
rect -722 -304 -721 -292
rect -974 -370 -973 -350
rect -971 -370 -970 -350
rect 272 -446 273 -406
rect 275 -446 276 -406
rect 342 -441 343 -421
rect 345 -441 346 -421
rect 385 -447 386 -407
rect 388 -447 389 -407
rect 614 -418 615 -393
rect 617 -418 618 -393
rect 622 -418 623 -393
rect 625 -418 626 -393
rect 652 -418 653 -393
rect 655 -418 656 -393
rect 696 -418 697 -393
rect 699 -418 700 -393
rect 741 -418 742 -393
rect 744 -418 745 -393
rect 309 -474 310 -454
rect 312 -474 313 -454
rect -1442 -606 -1441 -581
rect -1439 -606 -1438 -581
rect -1434 -606 -1433 -581
rect -1431 -606 -1430 -581
rect -1404 -606 -1403 -581
rect -1401 -606 -1400 -581
rect -1360 -606 -1359 -581
rect -1357 -606 -1356 -581
rect -1315 -606 -1314 -581
rect -1312 -606 -1311 -581
rect -1229 -606 -1228 -581
rect -1226 -606 -1225 -581
rect -1221 -606 -1220 -581
rect -1218 -606 -1217 -581
rect -1191 -606 -1190 -581
rect -1188 -606 -1187 -581
rect -1147 -606 -1146 -581
rect -1144 -606 -1143 -581
rect -1102 -606 -1101 -581
rect -1099 -606 -1098 -581
rect -982 -652 -981 -612
rect -979 -652 -978 -612
rect -736 -613 -735 -601
rect -733 -613 -731 -601
rect -727 -613 -725 -601
rect -723 -613 -722 -601
rect -912 -647 -911 -627
rect -909 -647 -908 -627
rect -869 -653 -868 -613
rect -866 -653 -865 -613
rect -696 -614 -695 -602
rect -693 -614 -692 -602
rect -945 -680 -944 -660
rect -942 -680 -941 -660
rect 293 -752 294 -712
rect 296 -752 297 -712
rect 363 -747 364 -727
rect 366 -747 367 -727
rect 406 -753 407 -713
rect 409 -753 410 -713
rect 635 -724 636 -699
rect 638 -724 639 -699
rect 643 -724 644 -699
rect 646 -724 647 -699
rect 673 -724 674 -699
rect 676 -724 677 -699
rect 717 -724 718 -699
rect 720 -724 721 -699
rect 762 -724 763 -699
rect 765 -724 766 -699
rect 330 -780 331 -760
rect 333 -780 334 -760
rect 700 -964 701 -939
rect 703 -964 704 -939
rect 708 -964 709 -939
rect 711 -964 712 -939
rect 738 -964 739 -939
rect 741 -964 742 -939
rect 782 -964 783 -939
rect 785 -964 786 -939
rect 827 -964 828 -939
rect 830 -964 831 -939
<< ndcontact >>
rect -1518 268 -1514 278
rect -1510 268 -1506 278
rect -1482 268 -1478 278
rect -1474 268 -1470 278
rect -1466 268 -1462 278
rect -1438 268 -1434 278
rect -1430 268 -1426 278
rect -1422 268 -1418 278
rect -1387 268 -1383 278
rect -1379 268 -1375 278
rect -1305 268 -1301 278
rect -1297 268 -1293 278
rect -1269 268 -1265 278
rect -1261 268 -1257 278
rect -1253 268 -1249 278
rect -1225 268 -1221 278
rect -1217 268 -1213 278
rect -1209 268 -1205 278
rect -1174 268 -1170 278
rect -1166 268 -1162 278
rect -1017 266 -1013 286
rect -1009 266 -1005 286
rect -808 261 -804 273
rect -790 261 -786 273
rect -768 272 -764 278
rect -760 272 -756 278
rect -1054 214 -1050 234
rect -1046 214 -1042 234
rect -984 219 -980 239
rect -976 219 -972 239
rect -941 213 -937 233
rect -933 213 -929 233
rect -629 230 -625 240
rect -621 230 -617 240
rect -593 230 -589 240
rect -585 230 -581 240
rect -577 230 -573 240
rect -549 230 -545 240
rect -541 230 -537 240
rect -533 230 -529 240
rect -498 230 -494 240
rect -490 230 -486 240
rect -115 149 -111 169
rect -107 149 -103 169
rect -77 149 -73 169
rect -69 149 -65 169
rect -33 149 -29 169
rect -25 149 -21 169
rect 5 149 9 169
rect 13 149 17 169
rect 291 133 295 153
rect 299 133 303 153
rect -158 11 -154 111
rect -150 11 -146 111
rect -80 10 -76 110
rect -72 10 -68 110
rect 254 81 258 101
rect 262 81 266 101
rect 324 86 328 106
rect 332 86 336 106
rect 592 117 596 127
rect 600 117 604 127
rect 628 117 632 127
rect 636 117 640 127
rect 644 117 648 127
rect 672 117 676 127
rect 680 117 684 127
rect 688 117 692 127
rect 723 117 727 127
rect 731 117 735 127
rect 367 80 371 100
rect 375 80 379 100
rect -1503 -61 -1499 -51
rect -1495 -61 -1491 -51
rect -1467 -61 -1463 -51
rect -1459 -61 -1455 -51
rect -1451 -61 -1447 -51
rect -1423 -61 -1419 -51
rect -1415 -61 -1411 -51
rect -1407 -61 -1403 -51
rect -1372 -61 -1368 -51
rect -1364 -61 -1360 -51
rect -1290 -61 -1286 -51
rect -1282 -61 -1278 -51
rect -1254 -61 -1250 -51
rect -1246 -61 -1242 -51
rect -1238 -61 -1234 -51
rect -1210 -61 -1206 -51
rect -1202 -61 -1198 -51
rect -1194 -61 -1190 -51
rect -1159 -61 -1155 -51
rect -1151 -61 -1147 -51
rect -1002 -63 -998 -43
rect -994 -63 -990 -43
rect -591 -50 -587 -44
rect -583 -50 -579 -44
rect -793 -68 -789 -56
rect -775 -68 -771 -56
rect -753 -57 -749 -51
rect -745 -57 -741 -51
rect -1039 -115 -1035 -95
rect -1031 -115 -1027 -95
rect -969 -110 -965 -90
rect -961 -110 -957 -90
rect -926 -116 -922 -96
rect -918 -116 -914 -96
rect -213 -127 -209 -27
rect -205 -127 -201 -27
rect -150 -128 -146 -28
rect -142 -128 -138 -28
rect -276 -272 -272 -172
rect -268 -272 -264 -172
rect -205 -272 -201 -172
rect -197 -272 -193 -172
rect 281 -175 285 -155
rect 289 -175 293 -155
rect 244 -227 248 -207
rect 252 -227 256 -207
rect 314 -222 318 -202
rect 322 -222 326 -202
rect 582 -191 586 -181
rect 590 -191 594 -181
rect 618 -191 622 -181
rect 626 -191 630 -181
rect 634 -191 638 -181
rect 662 -191 666 -181
rect 670 -191 674 -181
rect 678 -191 682 -181
rect 713 -191 717 -181
rect 721 -191 725 -181
rect 357 -228 361 -208
rect 365 -228 369 -208
rect -1479 -328 -1475 -318
rect -1471 -328 -1467 -318
rect -1443 -328 -1439 -318
rect -1435 -328 -1431 -318
rect -1427 -328 -1423 -318
rect -1399 -328 -1395 -318
rect -1391 -328 -1387 -318
rect -1383 -328 -1379 -318
rect -1348 -328 -1344 -318
rect -1340 -328 -1336 -318
rect -1266 -328 -1262 -318
rect -1258 -328 -1254 -318
rect -1230 -328 -1226 -318
rect -1222 -328 -1218 -318
rect -1214 -328 -1210 -318
rect -1186 -328 -1182 -318
rect -1178 -328 -1174 -318
rect -1170 -328 -1166 -318
rect -1135 -328 -1131 -318
rect -1127 -328 -1123 -318
rect -978 -330 -974 -310
rect -970 -330 -966 -310
rect -769 -335 -765 -323
rect -751 -335 -747 -323
rect -729 -324 -725 -318
rect -721 -324 -717 -318
rect -1015 -382 -1011 -362
rect -1007 -382 -1003 -362
rect -945 -377 -941 -357
rect -937 -377 -933 -357
rect -902 -383 -898 -363
rect -894 -383 -890 -363
rect -365 -420 -361 -320
rect -357 -420 -353 -320
rect -268 -420 -264 -320
rect -260 -420 -256 -320
rect 305 -434 309 -414
rect 313 -434 317 -414
rect -357 -565 -353 -465
rect -349 -565 -345 -465
rect 268 -486 272 -466
rect 276 -486 280 -466
rect 338 -481 342 -461
rect 346 -481 350 -461
rect 606 -450 610 -440
rect 614 -450 618 -440
rect 642 -450 646 -440
rect 650 -450 654 -440
rect 658 -450 662 -440
rect 686 -450 690 -440
rect 694 -450 698 -440
rect 702 -450 706 -440
rect 737 -450 741 -440
rect 745 -450 749 -440
rect 381 -487 385 -467
rect 389 -487 393 -467
rect -1450 -638 -1446 -628
rect -1442 -638 -1438 -628
rect -1414 -638 -1410 -628
rect -1406 -638 -1402 -628
rect -1398 -638 -1394 -628
rect -1370 -638 -1366 -628
rect -1362 -638 -1358 -628
rect -1354 -638 -1350 -628
rect -1319 -638 -1315 -628
rect -1311 -638 -1307 -628
rect -1237 -638 -1233 -628
rect -1229 -638 -1225 -628
rect -1201 -638 -1197 -628
rect -1193 -638 -1189 -628
rect -1185 -638 -1181 -628
rect -1157 -638 -1153 -628
rect -1149 -638 -1145 -628
rect -1141 -638 -1137 -628
rect -1106 -638 -1102 -628
rect -1098 -638 -1094 -628
rect -949 -640 -945 -620
rect -941 -640 -937 -620
rect -740 -645 -736 -633
rect -722 -645 -718 -633
rect -700 -634 -696 -628
rect -692 -634 -688 -628
rect -986 -692 -982 -672
rect -978 -692 -974 -672
rect -916 -687 -912 -667
rect -908 -687 -904 -667
rect -873 -693 -869 -673
rect -865 -693 -861 -673
rect -349 -698 -345 -598
rect -341 -698 -337 -598
rect 326 -740 330 -720
rect 334 -740 338 -720
rect 289 -792 293 -772
rect 297 -792 301 -772
rect 359 -787 363 -767
rect 367 -787 371 -767
rect 627 -756 631 -746
rect 635 -756 639 -746
rect 663 -756 667 -746
rect 671 -756 675 -746
rect 679 -756 683 -746
rect 707 -756 711 -746
rect 715 -756 719 -746
rect 723 -756 727 -746
rect 758 -756 762 -746
rect 766 -756 770 -746
rect 402 -793 406 -773
rect 410 -793 414 -773
rect 692 -996 696 -986
rect 700 -996 704 -986
rect 728 -996 732 -986
rect 736 -996 740 -986
rect 744 -996 748 -986
rect 772 -996 776 -986
rect 780 -996 784 -986
rect 788 -996 792 -986
rect 823 -996 827 -986
rect 831 -996 835 -986
<< pdcontact >>
rect -1514 300 -1510 325
rect -1506 300 -1502 325
rect -1498 300 -1494 325
rect -1476 300 -1472 325
rect -1468 300 -1464 325
rect -1432 300 -1428 325
rect -1424 300 -1420 325
rect -1387 300 -1383 325
rect -1379 300 -1375 325
rect -1301 300 -1297 325
rect -1293 300 -1289 325
rect -1285 300 -1281 325
rect -1263 300 -1259 325
rect -1255 300 -1251 325
rect -1219 300 -1215 325
rect -1211 300 -1207 325
rect -1174 300 -1170 325
rect -1166 300 -1162 325
rect -1054 254 -1050 294
rect -1046 254 -1042 294
rect -808 293 -804 305
rect -799 293 -795 305
rect -790 293 -786 305
rect -984 259 -980 279
rect -976 259 -972 279
rect -941 253 -937 293
rect -933 253 -929 293
rect -768 292 -764 304
rect -760 292 -756 304
rect -625 262 -621 287
rect -617 262 -613 287
rect -609 262 -605 287
rect -587 262 -583 287
rect -579 262 -575 287
rect -543 262 -539 287
rect -535 262 -531 287
rect -498 262 -494 287
rect -490 262 -486 287
rect -1017 226 -1013 246
rect -1009 226 -1005 246
rect -373 150 -369 200
rect -365 150 -361 200
rect -284 150 -280 200
rect -276 150 -272 200
rect -221 150 -217 200
rect -213 150 -209 200
rect -166 150 -162 200
rect -158 150 -154 200
rect -115 187 -111 227
rect -107 187 -103 227
rect -77 187 -73 227
rect -69 187 -65 227
rect -33 187 -29 227
rect -25 187 -21 227
rect 5 187 9 227
rect 13 187 17 227
rect 254 121 258 161
rect 262 121 266 161
rect 324 126 328 146
rect 332 126 336 146
rect 367 120 371 160
rect 375 120 379 160
rect 596 149 600 174
rect 604 149 608 174
rect 612 149 616 174
rect 634 149 638 174
rect 642 149 646 174
rect 678 149 682 174
rect 686 149 690 174
rect 723 149 727 174
rect 731 149 735 174
rect 291 93 295 113
rect 299 93 303 113
rect -1499 -29 -1495 -4
rect -1491 -29 -1487 -4
rect -1483 -29 -1479 -4
rect -1461 -29 -1457 -4
rect -1453 -29 -1449 -4
rect -1417 -29 -1413 -4
rect -1409 -29 -1405 -4
rect -1372 -29 -1368 -4
rect -1364 -29 -1360 -4
rect -1286 -29 -1282 -4
rect -1278 -29 -1274 -4
rect -1270 -29 -1266 -4
rect -1248 -29 -1244 -4
rect -1240 -29 -1236 -4
rect -1204 -29 -1200 -4
rect -1196 -29 -1192 -4
rect -1159 -29 -1155 -4
rect -1151 -29 -1147 -4
rect -1039 -75 -1035 -35
rect -1031 -75 -1027 -35
rect -793 -36 -789 -24
rect -784 -36 -780 -24
rect -775 -36 -771 -24
rect -969 -70 -965 -50
rect -961 -70 -957 -50
rect -926 -76 -922 -36
rect -918 -76 -914 -36
rect -753 -37 -749 -25
rect -745 -37 -741 -25
rect -591 -30 -587 -18
rect -583 -30 -579 -18
rect -1002 -103 -998 -83
rect -994 -103 -990 -83
rect -1475 -296 -1471 -271
rect -1467 -296 -1463 -271
rect -1459 -296 -1455 -271
rect -1437 -296 -1433 -271
rect -1429 -296 -1425 -271
rect -1393 -296 -1389 -271
rect -1385 -296 -1381 -271
rect -1348 -296 -1344 -271
rect -1340 -296 -1336 -271
rect -1262 -296 -1258 -271
rect -1254 -296 -1250 -271
rect -1246 -296 -1242 -271
rect -1224 -296 -1220 -271
rect -1216 -296 -1212 -271
rect -1180 -296 -1176 -271
rect -1172 -296 -1168 -271
rect -1135 -296 -1131 -271
rect -1127 -296 -1123 -271
rect 244 -187 248 -147
rect 252 -187 256 -147
rect 314 -182 318 -162
rect 322 -182 326 -162
rect 357 -188 361 -148
rect 365 -188 369 -148
rect 586 -159 590 -134
rect 594 -159 598 -134
rect 602 -159 606 -134
rect 624 -159 628 -134
rect 632 -159 636 -134
rect 668 -159 672 -134
rect 676 -159 680 -134
rect 713 -159 717 -134
rect 721 -159 725 -134
rect 281 -215 285 -195
rect 289 -215 293 -195
rect -1015 -342 -1011 -302
rect -1007 -342 -1003 -302
rect -769 -303 -765 -291
rect -760 -303 -756 -291
rect -751 -303 -747 -291
rect -945 -337 -941 -317
rect -937 -337 -933 -317
rect -902 -343 -898 -303
rect -894 -343 -890 -303
rect -729 -304 -725 -292
rect -721 -304 -717 -292
rect -978 -370 -974 -350
rect -970 -370 -966 -350
rect 268 -446 272 -406
rect 276 -446 280 -406
rect 338 -441 342 -421
rect 346 -441 350 -421
rect 381 -447 385 -407
rect 389 -447 393 -407
rect 610 -418 614 -393
rect 618 -418 622 -393
rect 626 -418 630 -393
rect 648 -418 652 -393
rect 656 -418 660 -393
rect 692 -418 696 -393
rect 700 -418 704 -393
rect 737 -418 741 -393
rect 745 -418 749 -393
rect 305 -474 309 -454
rect 313 -474 317 -454
rect -1446 -606 -1442 -581
rect -1438 -606 -1434 -581
rect -1430 -606 -1426 -581
rect -1408 -606 -1404 -581
rect -1400 -606 -1396 -581
rect -1364 -606 -1360 -581
rect -1356 -606 -1352 -581
rect -1319 -606 -1315 -581
rect -1311 -606 -1307 -581
rect -1233 -606 -1229 -581
rect -1225 -606 -1221 -581
rect -1217 -606 -1213 -581
rect -1195 -606 -1191 -581
rect -1187 -606 -1183 -581
rect -1151 -606 -1147 -581
rect -1143 -606 -1139 -581
rect -1106 -606 -1102 -581
rect -1098 -606 -1094 -581
rect -986 -652 -982 -612
rect -978 -652 -974 -612
rect -740 -613 -736 -601
rect -731 -613 -727 -601
rect -722 -613 -718 -601
rect -916 -647 -912 -627
rect -908 -647 -904 -627
rect -873 -653 -869 -613
rect -865 -653 -861 -613
rect -700 -614 -696 -602
rect -692 -614 -688 -602
rect -949 -680 -945 -660
rect -941 -680 -937 -660
rect 289 -752 293 -712
rect 297 -752 301 -712
rect 359 -747 363 -727
rect 367 -747 371 -727
rect 402 -753 406 -713
rect 410 -753 414 -713
rect 631 -724 635 -699
rect 639 -724 643 -699
rect 647 -724 651 -699
rect 669 -724 673 -699
rect 677 -724 681 -699
rect 713 -724 717 -699
rect 721 -724 725 -699
rect 758 -724 762 -699
rect 766 -724 770 -699
rect 326 -780 330 -760
rect 334 -780 338 -760
rect 696 -964 700 -939
rect 704 -964 708 -939
rect 712 -964 716 -939
rect 734 -964 738 -939
rect 742 -964 746 -939
rect 778 -964 782 -939
rect 786 -964 790 -939
rect 823 -964 827 -939
rect 831 -964 835 -939
<< nsubstratencontact >>
rect -120 233 -116 237
rect -82 233 -78 237
rect -38 233 -34 237
rect 0 233 4 237
rect -378 206 -374 210
rect -289 206 -285 210
rect -226 206 -222 210
rect -171 206 -167 210
<< polysilicon >>
rect -1509 325 -1507 328
rect -1501 325 -1499 328
rect -1471 325 -1469 328
rect -1427 325 -1425 328
rect -1382 325 -1380 328
rect -1296 325 -1294 328
rect -1288 325 -1286 328
rect -1258 325 -1256 328
rect -1214 325 -1212 328
rect -1169 325 -1167 328
rect -803 305 -801 308
rect -793 305 -791 308
rect -1509 293 -1507 300
rect -1514 289 -1507 293
rect -1513 278 -1511 289
rect -1501 281 -1499 300
rect -1471 292 -1469 300
rect -1427 292 -1425 300
rect -1477 290 -1469 292
rect -1433 290 -1425 292
rect -1477 278 -1475 290
rect -1469 278 -1467 287
rect -1433 278 -1431 290
rect -1425 278 -1423 287
rect -1382 278 -1380 300
rect -1296 293 -1294 300
rect -1301 289 -1294 293
rect -1300 278 -1298 289
rect -1288 281 -1286 300
rect -1258 292 -1256 300
rect -1214 292 -1212 300
rect -1264 290 -1256 292
rect -1220 290 -1212 292
rect -1264 278 -1262 290
rect -1256 278 -1254 287
rect -1220 278 -1218 290
rect -1212 278 -1210 287
rect -1169 278 -1167 300
rect -1049 294 -1047 298
rect -1513 265 -1511 268
rect -1477 265 -1475 268
rect -1469 265 -1467 268
rect -1433 265 -1431 268
rect -1425 265 -1423 268
rect -1382 265 -1380 268
rect -1300 265 -1298 268
rect -1264 265 -1262 268
rect -1256 265 -1254 268
rect -1220 265 -1218 268
rect -1212 265 -1210 268
rect -1169 265 -1167 268
rect -936 293 -934 297
rect -763 304 -761 307
rect -1012 286 -1010 293
rect -979 279 -977 293
rect -1012 263 -1010 266
rect -979 256 -977 259
rect -1049 234 -1047 254
rect -803 273 -801 293
rect -793 273 -791 293
rect -763 278 -761 292
rect -620 287 -618 290
rect -612 287 -610 290
rect -582 287 -580 290
rect -538 287 -536 290
rect -493 287 -491 290
rect -763 269 -761 272
rect -803 258 -801 261
rect -793 258 -791 261
rect -620 255 -618 262
rect -1012 246 -1010 249
rect -979 239 -977 242
rect -1049 211 -1047 214
rect -1012 212 -1010 226
rect -936 233 -934 253
rect -625 251 -618 255
rect -624 240 -622 251
rect -612 243 -610 262
rect -582 254 -580 262
rect -538 254 -536 262
rect -588 252 -580 254
rect -544 252 -536 254
rect -588 240 -586 252
rect -580 240 -578 249
rect -544 240 -542 252
rect -536 240 -534 249
rect -493 240 -491 262
rect -979 212 -977 219
rect -624 227 -622 230
rect -588 227 -586 230
rect -580 227 -578 230
rect -544 227 -542 230
rect -536 227 -534 230
rect -493 227 -491 230
rect -110 227 -108 230
rect -72 227 -70 230
rect -28 227 -26 230
rect 10 227 12 230
rect -936 210 -934 213
rect -368 200 -366 203
rect -279 200 -277 203
rect -216 200 -214 203
rect -161 200 -159 203
rect -110 169 -108 187
rect -72 169 -70 187
rect -28 169 -26 187
rect 10 169 12 187
rect 601 174 603 177
rect 609 174 611 177
rect 639 174 641 177
rect 683 174 685 177
rect 728 174 730 177
rect -368 133 -366 150
rect -279 133 -277 150
rect -216 133 -214 150
rect -161 133 -159 150
rect 259 161 261 165
rect -110 145 -108 149
rect -72 145 -70 149
rect -28 145 -26 149
rect 10 145 12 149
rect 372 160 374 164
rect 296 153 298 160
rect 329 146 331 160
rect 296 130 298 133
rect 329 123 331 126
rect -153 111 -151 114
rect -75 110 -73 113
rect -153 -1 -151 11
rect 259 101 261 121
rect 601 142 603 149
rect 596 138 603 142
rect 597 127 599 138
rect 609 130 611 149
rect 639 141 641 149
rect 683 141 685 149
rect 633 139 641 141
rect 677 139 685 141
rect 633 127 635 139
rect 641 127 643 136
rect 677 127 679 139
rect 685 127 687 136
rect 728 127 730 149
rect 296 113 298 116
rect 329 106 331 109
rect 259 78 261 81
rect 296 79 298 93
rect 372 100 374 120
rect 597 114 599 117
rect 633 114 635 117
rect 641 114 643 117
rect 677 114 679 117
rect 685 114 687 117
rect 728 114 730 117
rect 329 79 331 86
rect 372 77 374 80
rect -1494 -4 -1492 -1
rect -1486 -4 -1484 -1
rect -1456 -4 -1454 -1
rect -1412 -4 -1410 -1
rect -1367 -4 -1365 -1
rect -1281 -4 -1279 -1
rect -1273 -4 -1271 -1
rect -1243 -4 -1241 -1
rect -1199 -4 -1197 -1
rect -1154 -4 -1152 -1
rect -75 -2 -73 10
rect -586 -18 -584 -15
rect -788 -24 -786 -21
rect -778 -24 -776 -21
rect -1494 -36 -1492 -29
rect -1499 -40 -1492 -36
rect -1498 -51 -1496 -40
rect -1486 -48 -1484 -29
rect -1456 -37 -1454 -29
rect -1412 -37 -1410 -29
rect -1462 -39 -1454 -37
rect -1418 -39 -1410 -37
rect -1462 -51 -1460 -39
rect -1454 -51 -1452 -42
rect -1418 -51 -1416 -39
rect -1410 -51 -1408 -42
rect -1367 -51 -1365 -29
rect -1281 -36 -1279 -29
rect -1286 -40 -1279 -36
rect -1285 -51 -1283 -40
rect -1273 -48 -1271 -29
rect -1243 -37 -1241 -29
rect -1199 -37 -1197 -29
rect -1249 -39 -1241 -37
rect -1205 -39 -1197 -37
rect -1249 -51 -1247 -39
rect -1241 -51 -1239 -42
rect -1205 -51 -1203 -39
rect -1197 -51 -1195 -42
rect -1154 -51 -1152 -29
rect -1034 -35 -1032 -31
rect -1498 -64 -1496 -61
rect -1462 -64 -1460 -61
rect -1454 -64 -1452 -61
rect -1418 -64 -1416 -61
rect -1410 -64 -1408 -61
rect -1367 -64 -1365 -61
rect -1285 -64 -1283 -61
rect -1249 -64 -1247 -61
rect -1241 -64 -1239 -61
rect -1205 -64 -1203 -61
rect -1197 -64 -1195 -61
rect -1154 -64 -1152 -61
rect -921 -36 -919 -32
rect -748 -25 -746 -22
rect -997 -43 -995 -36
rect -964 -50 -962 -36
rect -997 -66 -995 -63
rect -964 -73 -962 -70
rect -1034 -95 -1032 -75
rect -788 -56 -786 -36
rect -778 -56 -776 -36
rect -208 -27 -206 -24
rect -748 -51 -746 -37
rect -586 -44 -584 -30
rect -586 -53 -584 -50
rect -748 -60 -746 -57
rect -788 -71 -786 -68
rect -778 -71 -776 -68
rect -997 -83 -995 -80
rect -964 -90 -962 -87
rect -1034 -118 -1032 -115
rect -997 -117 -995 -103
rect -921 -96 -919 -76
rect -964 -117 -962 -110
rect -921 -119 -919 -116
rect -145 -28 -143 -25
rect -208 -139 -206 -127
rect -145 -140 -143 -128
rect 591 -134 593 -131
rect 599 -134 601 -131
rect 629 -134 631 -131
rect 673 -134 675 -131
rect 718 -134 720 -131
rect 249 -147 251 -143
rect -271 -172 -269 -169
rect -200 -172 -198 -169
rect -1470 -271 -1468 -268
rect -1462 -271 -1460 -268
rect -1432 -271 -1430 -268
rect -1388 -271 -1386 -268
rect -1343 -271 -1341 -268
rect -1257 -271 -1255 -268
rect -1249 -271 -1247 -268
rect -1219 -271 -1217 -268
rect -1175 -271 -1173 -268
rect -1130 -271 -1128 -268
rect 362 -148 364 -144
rect 286 -155 288 -148
rect 319 -162 321 -148
rect 286 -178 288 -175
rect 319 -185 321 -182
rect 249 -207 251 -187
rect 591 -166 593 -159
rect 586 -170 593 -166
rect 587 -181 589 -170
rect 599 -178 601 -159
rect 629 -167 631 -159
rect 673 -167 675 -159
rect 623 -169 631 -167
rect 667 -169 675 -167
rect 623 -181 625 -169
rect 631 -181 633 -172
rect 667 -181 669 -169
rect 675 -181 677 -172
rect 718 -181 720 -159
rect 286 -195 288 -192
rect 319 -202 321 -199
rect 249 -230 251 -227
rect 286 -229 288 -215
rect 362 -208 364 -188
rect 587 -194 589 -191
rect 623 -194 625 -191
rect 631 -194 633 -191
rect 667 -194 669 -191
rect 675 -194 677 -191
rect 718 -194 720 -191
rect 319 -229 321 -222
rect 362 -231 364 -228
rect -271 -284 -269 -272
rect -200 -284 -198 -272
rect -764 -291 -762 -288
rect -754 -291 -752 -288
rect -1470 -303 -1468 -296
rect -1475 -307 -1468 -303
rect -1474 -318 -1472 -307
rect -1462 -315 -1460 -296
rect -1432 -304 -1430 -296
rect -1388 -304 -1386 -296
rect -1438 -306 -1430 -304
rect -1394 -306 -1386 -304
rect -1438 -318 -1436 -306
rect -1430 -318 -1428 -309
rect -1394 -318 -1392 -306
rect -1386 -318 -1384 -309
rect -1343 -318 -1341 -296
rect -1257 -303 -1255 -296
rect -1262 -307 -1255 -303
rect -1261 -318 -1259 -307
rect -1249 -315 -1247 -296
rect -1219 -304 -1217 -296
rect -1175 -304 -1173 -296
rect -1225 -306 -1217 -304
rect -1181 -306 -1173 -304
rect -1225 -318 -1223 -306
rect -1217 -318 -1215 -309
rect -1181 -318 -1179 -306
rect -1173 -318 -1171 -309
rect -1130 -318 -1128 -296
rect -1010 -302 -1008 -298
rect -1474 -331 -1472 -328
rect -1438 -331 -1436 -328
rect -1430 -331 -1428 -328
rect -1394 -331 -1392 -328
rect -1386 -331 -1384 -328
rect -1343 -331 -1341 -328
rect -1261 -331 -1259 -328
rect -1225 -331 -1223 -328
rect -1217 -331 -1215 -328
rect -1181 -331 -1179 -328
rect -1173 -331 -1171 -328
rect -1130 -331 -1128 -328
rect -897 -303 -895 -299
rect -724 -292 -722 -289
rect -973 -310 -971 -303
rect -940 -317 -938 -303
rect -973 -333 -971 -330
rect -940 -340 -938 -337
rect -1010 -362 -1008 -342
rect -764 -323 -762 -303
rect -754 -323 -752 -303
rect -724 -318 -722 -304
rect -360 -320 -358 -317
rect -263 -320 -261 -317
rect -724 -327 -722 -324
rect -764 -338 -762 -335
rect -754 -338 -752 -335
rect -973 -350 -971 -347
rect -940 -357 -938 -354
rect -1010 -385 -1008 -382
rect -973 -384 -971 -370
rect -897 -363 -895 -343
rect -940 -384 -938 -377
rect -897 -386 -895 -383
rect 615 -393 617 -390
rect 623 -393 625 -390
rect 653 -393 655 -390
rect 697 -393 699 -390
rect 742 -393 744 -390
rect 273 -406 275 -402
rect -360 -432 -358 -420
rect -263 -432 -261 -420
rect 386 -407 388 -403
rect 310 -414 312 -407
rect 343 -421 345 -407
rect 310 -437 312 -434
rect 343 -444 345 -441
rect -352 -465 -350 -462
rect 273 -466 275 -446
rect 615 -425 617 -418
rect 610 -429 617 -425
rect 611 -440 613 -429
rect 623 -437 625 -418
rect 653 -426 655 -418
rect 697 -426 699 -418
rect 647 -428 655 -426
rect 691 -428 699 -426
rect 647 -440 649 -428
rect 655 -440 657 -431
rect 691 -440 693 -428
rect 699 -440 701 -431
rect 742 -440 744 -418
rect 310 -454 312 -451
rect 343 -461 345 -458
rect 273 -489 275 -486
rect 310 -488 312 -474
rect 386 -467 388 -447
rect 611 -453 613 -450
rect 647 -453 649 -450
rect 655 -453 657 -450
rect 691 -453 693 -450
rect 699 -453 701 -450
rect 742 -453 744 -450
rect 343 -488 345 -481
rect 386 -490 388 -487
rect -352 -577 -350 -565
rect -1441 -581 -1439 -578
rect -1433 -581 -1431 -578
rect -1403 -581 -1401 -578
rect -1359 -581 -1357 -578
rect -1314 -581 -1312 -578
rect -1228 -581 -1226 -578
rect -1220 -581 -1218 -578
rect -1190 -581 -1188 -578
rect -1146 -581 -1144 -578
rect -1101 -581 -1099 -578
rect -344 -598 -342 -595
rect -735 -601 -733 -598
rect -725 -601 -723 -598
rect -1441 -613 -1439 -606
rect -1446 -617 -1439 -613
rect -1445 -628 -1443 -617
rect -1433 -625 -1431 -606
rect -1403 -614 -1401 -606
rect -1359 -614 -1357 -606
rect -1409 -616 -1401 -614
rect -1365 -616 -1357 -614
rect -1409 -628 -1407 -616
rect -1401 -628 -1399 -619
rect -1365 -628 -1363 -616
rect -1357 -628 -1355 -619
rect -1314 -628 -1312 -606
rect -1228 -613 -1226 -606
rect -1233 -617 -1226 -613
rect -1232 -628 -1230 -617
rect -1220 -625 -1218 -606
rect -1190 -614 -1188 -606
rect -1146 -614 -1144 -606
rect -1196 -616 -1188 -614
rect -1152 -616 -1144 -614
rect -1196 -628 -1194 -616
rect -1188 -628 -1186 -619
rect -1152 -628 -1150 -616
rect -1144 -628 -1142 -619
rect -1101 -628 -1099 -606
rect -981 -612 -979 -608
rect -1445 -641 -1443 -638
rect -1409 -641 -1407 -638
rect -1401 -641 -1399 -638
rect -1365 -641 -1363 -638
rect -1357 -641 -1355 -638
rect -1314 -641 -1312 -638
rect -1232 -641 -1230 -638
rect -1196 -641 -1194 -638
rect -1188 -641 -1186 -638
rect -1152 -641 -1150 -638
rect -1144 -641 -1142 -638
rect -1101 -641 -1099 -638
rect -868 -613 -866 -609
rect -695 -602 -693 -599
rect -944 -620 -942 -613
rect -911 -627 -909 -613
rect -944 -643 -942 -640
rect -911 -650 -909 -647
rect -981 -672 -979 -652
rect -735 -633 -733 -613
rect -725 -633 -723 -613
rect -695 -628 -693 -614
rect -695 -637 -693 -634
rect -735 -648 -733 -645
rect -725 -648 -723 -645
rect -944 -660 -942 -657
rect -911 -667 -909 -664
rect -981 -695 -979 -692
rect -944 -694 -942 -680
rect -868 -673 -866 -653
rect -911 -694 -909 -687
rect -868 -696 -866 -693
rect -344 -710 -342 -698
rect 636 -699 638 -696
rect 644 -699 646 -696
rect 674 -699 676 -696
rect 718 -699 720 -696
rect 763 -699 765 -696
rect 294 -712 296 -708
rect 407 -713 409 -709
rect 331 -720 333 -713
rect 364 -727 366 -713
rect 331 -743 333 -740
rect 364 -750 366 -747
rect 294 -772 296 -752
rect 636 -731 638 -724
rect 631 -735 638 -731
rect 632 -746 634 -735
rect 644 -743 646 -724
rect 674 -732 676 -724
rect 718 -732 720 -724
rect 668 -734 676 -732
rect 712 -734 720 -732
rect 668 -746 670 -734
rect 676 -746 678 -737
rect 712 -746 714 -734
rect 720 -746 722 -737
rect 763 -746 765 -724
rect 331 -760 333 -757
rect 364 -767 366 -764
rect 294 -795 296 -792
rect 331 -794 333 -780
rect 407 -773 409 -753
rect 632 -759 634 -756
rect 668 -759 670 -756
rect 676 -759 678 -756
rect 712 -759 714 -756
rect 720 -759 722 -756
rect 763 -759 765 -756
rect 364 -794 366 -787
rect 407 -796 409 -793
rect 701 -939 703 -936
rect 709 -939 711 -936
rect 739 -939 741 -936
rect 783 -939 785 -936
rect 828 -939 830 -936
rect 701 -971 703 -964
rect 696 -975 703 -971
rect 697 -986 699 -975
rect 709 -983 711 -964
rect 739 -972 741 -964
rect 783 -972 785 -964
rect 733 -974 741 -972
rect 777 -974 785 -972
rect 733 -986 735 -974
rect 741 -986 743 -977
rect 777 -986 779 -974
rect 785 -986 787 -977
rect 828 -986 830 -964
rect 697 -999 699 -996
rect 733 -999 735 -996
rect 741 -999 743 -996
rect 777 -999 779 -996
rect 785 -999 787 -996
rect 828 -999 830 -996
<< polycontact >>
rect -1518 289 -1514 293
rect -1505 281 -1501 285
rect -1482 281 -1477 286
rect -1467 281 -1462 285
rect -1438 281 -1433 286
rect -1386 286 -1382 291
rect -1423 281 -1418 285
rect -1305 289 -1301 293
rect -1292 281 -1288 285
rect -1269 281 -1264 286
rect -1254 281 -1249 285
rect -1225 281 -1220 286
rect -1173 286 -1169 291
rect -1210 281 -1205 285
rect -1013 293 -1009 298
rect -980 293 -976 298
rect -1053 237 -1049 242
rect -807 282 -803 286
rect -797 276 -793 280
rect -767 281 -763 285
rect -940 236 -936 241
rect -629 251 -625 255
rect -616 243 -612 247
rect -593 243 -588 248
rect -578 243 -573 247
rect -549 243 -544 248
rect -497 248 -493 253
rect -534 243 -529 247
rect -1013 207 -1009 212
rect -980 207 -976 212
rect 295 160 299 165
rect 328 160 332 165
rect 255 104 259 109
rect 592 138 596 142
rect 605 130 609 134
rect 628 130 633 135
rect 643 130 648 134
rect 672 130 677 135
rect 724 135 728 140
rect 687 130 692 134
rect 368 103 372 108
rect 295 74 299 79
rect 328 74 332 79
rect -1503 -40 -1499 -36
rect -1490 -48 -1486 -44
rect -1467 -48 -1462 -43
rect -1452 -48 -1447 -44
rect -1423 -48 -1418 -43
rect -1371 -43 -1367 -38
rect -1408 -48 -1403 -44
rect -1290 -40 -1286 -36
rect -1277 -48 -1273 -44
rect -1254 -48 -1249 -43
rect -1239 -48 -1234 -44
rect -1210 -48 -1205 -43
rect -1158 -43 -1154 -38
rect -1195 -48 -1190 -44
rect -998 -36 -994 -31
rect -965 -36 -961 -31
rect -1038 -92 -1034 -87
rect -792 -47 -788 -43
rect -782 -53 -778 -49
rect -752 -48 -748 -44
rect -590 -41 -586 -37
rect -925 -93 -921 -88
rect -998 -122 -994 -117
rect -965 -122 -961 -117
rect 285 -148 289 -143
rect 318 -148 322 -143
rect 245 -204 249 -199
rect 582 -170 586 -166
rect 595 -178 599 -174
rect 618 -178 623 -173
rect 633 -178 638 -174
rect 662 -178 667 -173
rect 714 -173 718 -168
rect 677 -178 682 -174
rect 358 -205 362 -200
rect 285 -234 289 -229
rect 318 -234 322 -229
rect -1479 -307 -1475 -303
rect -1466 -315 -1462 -311
rect -1443 -315 -1438 -310
rect -1428 -315 -1423 -311
rect -1399 -315 -1394 -310
rect -1347 -310 -1343 -305
rect -1384 -315 -1379 -311
rect -1266 -307 -1262 -303
rect -1253 -315 -1249 -311
rect -1230 -315 -1225 -310
rect -1215 -315 -1210 -311
rect -1186 -315 -1181 -310
rect -1134 -310 -1130 -305
rect -1171 -315 -1166 -311
rect -974 -303 -970 -298
rect -941 -303 -937 -298
rect -1014 -359 -1010 -354
rect -768 -314 -764 -310
rect -758 -320 -754 -316
rect -728 -315 -724 -311
rect -901 -360 -897 -355
rect -974 -389 -970 -384
rect -941 -389 -937 -384
rect 309 -407 313 -402
rect 342 -407 346 -402
rect 269 -463 273 -458
rect 606 -429 610 -425
rect 619 -437 623 -433
rect 642 -437 647 -432
rect 657 -437 662 -433
rect 686 -437 691 -432
rect 738 -432 742 -427
rect 701 -437 706 -433
rect 382 -464 386 -459
rect 309 -493 313 -488
rect 342 -493 346 -488
rect -1450 -617 -1446 -613
rect -1437 -625 -1433 -621
rect -1414 -625 -1409 -620
rect -1399 -625 -1394 -621
rect -1370 -625 -1365 -620
rect -1318 -620 -1314 -615
rect -1355 -625 -1350 -621
rect -1237 -617 -1233 -613
rect -1224 -625 -1220 -621
rect -1201 -625 -1196 -620
rect -1186 -625 -1181 -621
rect -1157 -625 -1152 -620
rect -1105 -620 -1101 -615
rect -1142 -625 -1137 -621
rect -945 -613 -941 -608
rect -912 -613 -908 -608
rect -985 -669 -981 -664
rect -739 -624 -735 -620
rect -729 -630 -725 -626
rect -699 -625 -695 -621
rect -872 -670 -868 -665
rect -945 -699 -941 -694
rect -912 -699 -908 -694
rect 330 -713 334 -708
rect 363 -713 367 -708
rect 290 -769 294 -764
rect 627 -735 631 -731
rect 640 -743 644 -739
rect 663 -743 668 -738
rect 678 -743 683 -739
rect 707 -743 712 -738
rect 759 -738 763 -733
rect 722 -743 727 -739
rect 403 -770 407 -765
rect 330 -799 334 -794
rect 363 -799 367 -794
rect 692 -975 696 -971
rect 705 -983 709 -979
rect 728 -983 733 -978
rect 743 -983 748 -979
rect 772 -983 777 -978
rect 824 -978 828 -973
rect 787 -983 792 -979
<< metal1 >>
rect -1520 331 -816 335
rect -1514 325 -1510 331
rect -1476 325 -1472 331
rect -1432 325 -1428 331
rect -1387 325 -1383 331
rect -1301 325 -1297 331
rect -1263 325 -1259 331
rect -1219 325 -1215 331
rect -1174 325 -1170 331
rect -1082 330 -816 331
rect -1464 300 -1451 325
rect -1420 300 -1407 325
rect -1251 300 -1238 325
rect -1207 300 -1194 325
rect -1525 289 -1518 293
rect -1498 292 -1494 300
rect -1498 289 -1458 292
rect -1508 281 -1505 285
rect -1498 278 -1494 289
rect -1486 281 -1482 286
rect -1462 281 -1458 289
rect -1454 286 -1451 300
rect -1410 291 -1407 300
rect -1410 286 -1386 291
rect -1379 290 -1375 300
rect -1454 281 -1438 286
rect -1418 281 -1414 285
rect -1454 278 -1451 281
rect -1410 278 -1407 286
rect -1379 285 -1366 290
rect -1379 278 -1375 285
rect -1312 289 -1305 293
rect -1285 292 -1281 300
rect -1285 289 -1245 292
rect -1295 281 -1292 285
rect -1285 278 -1281 289
rect -1273 281 -1269 286
rect -1249 281 -1245 289
rect -1241 286 -1238 300
rect -1197 291 -1194 300
rect -1197 286 -1173 291
rect -1166 290 -1162 300
rect -1054 294 -1050 330
rect -1241 281 -1225 286
rect -1205 281 -1201 285
rect -1241 278 -1238 281
rect -1197 278 -1194 286
rect -1166 285 -1153 290
rect -1166 278 -1162 285
rect -1506 268 -1494 278
rect -1462 268 -1451 278
rect -1418 268 -1407 278
rect -1293 268 -1281 278
rect -1249 268 -1238 278
rect -1205 268 -1194 278
rect -1518 263 -1514 268
rect -1482 263 -1478 268
rect -1438 263 -1434 268
rect -1387 263 -1383 268
rect -1305 263 -1301 268
rect -1269 263 -1265 268
rect -1225 263 -1221 268
rect -1174 263 -1170 268
rect -1519 259 -1162 263
rect -1166 174 -1162 259
rect -1029 262 -1024 317
rect -1013 298 -1009 305
rect -980 298 -976 305
rect -941 293 -937 330
rect -854 310 -848 317
rect -821 314 -816 330
rect -821 313 -771 314
rect -821 311 -750 313
rect -921 305 -840 310
rect -1017 262 -1013 266
rect -1029 258 -1013 262
rect -1063 237 -1053 242
rect -1046 241 -1042 254
rect -1017 246 -1013 258
rect -1046 236 -1033 241
rect -1046 234 -1042 236
rect -1009 261 -1005 266
rect -1009 257 -992 261
rect -1009 246 -1005 257
rect -996 247 -992 257
rect -984 247 -980 259
rect -996 242 -980 247
rect -1054 175 -1050 214
rect -1013 194 -1009 207
rect -996 181 -990 242
rect -984 239 -980 242
rect -976 246 -972 259
rect -976 242 -955 246
rect -976 239 -972 242
rect -961 241 -955 242
rect -961 236 -951 241
rect -945 236 -940 241
rect -933 240 -929 253
rect -891 279 -882 292
rect -843 285 -840 305
rect -808 305 -805 311
rect -789 305 -786 311
rect -774 310 -750 311
rect -768 304 -765 310
rect -799 290 -796 293
rect -631 293 -478 297
rect -799 287 -786 290
rect -843 282 -807 285
rect -789 284 -786 287
rect -789 281 -767 284
rect -759 284 -756 292
rect -625 287 -621 293
rect -587 287 -583 293
rect -543 287 -539 293
rect -498 287 -494 293
rect -759 281 -747 284
rect -891 276 -797 279
rect -933 235 -916 240
rect -933 233 -929 235
rect -980 194 -976 207
rect -941 175 -937 213
rect -891 195 -883 276
rect -789 273 -786 281
rect -759 278 -756 281
rect -768 268 -765 272
rect -778 265 -750 268
rect -808 255 -805 261
rect -778 255 -774 265
rect -575 262 -562 287
rect -531 262 -518 287
rect -873 252 -774 255
rect -873 175 -862 252
rect -636 251 -629 255
rect -609 254 -605 262
rect -609 251 -569 254
rect -619 243 -616 247
rect -609 240 -605 251
rect -597 243 -593 248
rect -573 243 -569 251
rect -565 248 -562 262
rect -521 253 -518 262
rect -521 248 -497 253
rect -490 252 -486 262
rect -565 243 -549 248
rect -529 243 -525 247
rect -565 240 -562 243
rect -521 240 -518 248
rect -490 247 -477 252
rect -490 240 -486 247
rect -121 240 23 245
rect -617 230 -605 240
rect -573 230 -562 240
rect -529 230 -518 240
rect -115 237 -111 240
rect -77 237 -73 240
rect -33 237 -29 240
rect 5 237 9 240
rect -121 233 -120 237
rect -116 233 -111 237
rect -83 233 -82 237
rect -78 233 -73 237
rect -39 233 -38 237
rect -34 233 -29 237
rect -1 233 0 237
rect 4 233 9 237
rect -629 225 -625 230
rect -593 225 -589 230
rect -549 225 -545 230
rect -498 225 -494 230
rect -115 227 -111 233
rect -77 227 -73 233
rect -33 227 -29 233
rect 5 227 9 233
rect -630 221 -486 225
rect -373 210 -369 219
rect -284 210 -280 219
rect -221 210 -217 219
rect -166 210 -162 219
rect -379 206 -378 210
rect -374 206 -369 210
rect -290 206 -289 210
rect -285 206 -280 210
rect -227 206 -226 210
rect -222 206 -217 210
rect -172 206 -171 210
rect -167 206 -162 210
rect -1082 174 -862 175
rect -1166 167 -862 174
rect -373 200 -369 206
rect -284 200 -280 206
rect -221 200 -217 206
rect -166 200 -162 206
rect 226 197 459 202
rect -107 169 -103 187
rect -69 169 -65 187
rect -25 169 -21 187
rect 13 169 17 187
rect -1505 2 -801 6
rect -1499 -4 -1495 2
rect -1461 -4 -1457 2
rect -1417 -4 -1413 2
rect -1372 -4 -1368 2
rect -1286 -4 -1282 2
rect -1248 -4 -1244 2
rect -1204 -4 -1200 2
rect -1159 -4 -1155 2
rect -1067 1 -801 2
rect -1449 -29 -1436 -4
rect -1405 -29 -1392 -4
rect -1236 -29 -1223 -4
rect -1192 -29 -1179 -4
rect -1510 -40 -1503 -36
rect -1483 -37 -1479 -29
rect -1483 -40 -1443 -37
rect -1493 -48 -1490 -44
rect -1483 -51 -1479 -40
rect -1471 -48 -1467 -43
rect -1447 -48 -1443 -40
rect -1439 -43 -1436 -29
rect -1395 -38 -1392 -29
rect -1395 -43 -1371 -38
rect -1364 -39 -1360 -29
rect -1439 -48 -1423 -43
rect -1403 -48 -1399 -44
rect -1439 -51 -1436 -48
rect -1395 -51 -1392 -43
rect -1364 -44 -1351 -39
rect -1364 -51 -1360 -44
rect -1297 -40 -1290 -36
rect -1270 -37 -1266 -29
rect -1270 -40 -1230 -37
rect -1280 -48 -1277 -44
rect -1270 -51 -1266 -40
rect -1258 -48 -1254 -43
rect -1234 -48 -1230 -40
rect -1226 -43 -1223 -29
rect -1182 -38 -1179 -29
rect -1182 -43 -1158 -38
rect -1151 -39 -1147 -29
rect -1039 -35 -1035 1
rect -1226 -48 -1210 -43
rect -1190 -48 -1186 -44
rect -1226 -51 -1223 -48
rect -1182 -51 -1179 -43
rect -1151 -44 -1138 -39
rect -1151 -51 -1147 -44
rect -1491 -61 -1479 -51
rect -1447 -61 -1436 -51
rect -1403 -61 -1392 -51
rect -1278 -61 -1266 -51
rect -1234 -61 -1223 -51
rect -1190 -61 -1179 -51
rect -1503 -66 -1499 -61
rect -1467 -66 -1463 -61
rect -1423 -66 -1419 -61
rect -1372 -66 -1368 -61
rect -1290 -66 -1286 -61
rect -1254 -66 -1250 -61
rect -1210 -66 -1206 -61
rect -1159 -66 -1155 -61
rect -1504 -70 -1147 -66
rect -1151 -155 -1147 -70
rect -1014 -67 -1009 -12
rect -998 -31 -994 -24
rect -965 -31 -961 -24
rect -926 -36 -922 1
rect -839 -19 -833 -12
rect -806 -15 -801 1
rect -597 -12 -573 -9
rect -806 -16 -756 -15
rect -806 -18 -735 -16
rect -906 -24 -825 -19
rect -1002 -67 -998 -63
rect -1014 -71 -998 -67
rect -1048 -92 -1038 -87
rect -1031 -88 -1027 -75
rect -1002 -83 -998 -71
rect -1031 -93 -1018 -88
rect -1031 -95 -1027 -93
rect -994 -68 -990 -63
rect -994 -72 -977 -68
rect -994 -83 -990 -72
rect -981 -82 -977 -72
rect -969 -82 -965 -70
rect -981 -87 -965 -82
rect -1039 -154 -1035 -115
rect -998 -135 -994 -122
rect -981 -148 -975 -87
rect -969 -90 -965 -87
rect -961 -83 -957 -70
rect -961 -87 -940 -83
rect -961 -90 -957 -87
rect -946 -88 -940 -87
rect -946 -93 -936 -88
rect -930 -93 -925 -88
rect -918 -89 -914 -76
rect -876 -50 -867 -37
rect -828 -44 -825 -24
rect -793 -24 -790 -18
rect -774 -24 -771 -18
rect -759 -19 -735 -18
rect -591 -18 -588 -12
rect -753 -25 -750 -19
rect -784 -39 -781 -36
rect -784 -42 -771 -39
rect -828 -47 -792 -44
rect -774 -45 -771 -42
rect -774 -48 -752 -45
rect -744 -45 -741 -37
rect -597 -41 -590 -38
rect -582 -38 -579 -30
rect -582 -41 -573 -38
rect -582 -44 -579 -41
rect -744 -48 -732 -45
rect -876 -53 -782 -50
rect -918 -94 -901 -89
rect -918 -96 -914 -94
rect -965 -135 -961 -122
rect -926 -154 -922 -116
rect -876 -134 -868 -53
rect -774 -56 -771 -48
rect -744 -51 -741 -48
rect -591 -54 -588 -50
rect -597 -57 -573 -54
rect -753 -61 -750 -57
rect -763 -64 -735 -61
rect -793 -74 -790 -68
rect -763 -74 -759 -64
rect -858 -77 -759 -74
rect -858 -154 -847 -77
rect -1067 -155 -847 -154
rect -1151 -162 -847 -155
rect -1481 -265 -777 -261
rect -1475 -271 -1471 -265
rect -1437 -271 -1433 -265
rect -1393 -271 -1389 -265
rect -1348 -271 -1344 -265
rect -1262 -271 -1258 -265
rect -1224 -271 -1220 -265
rect -1180 -271 -1176 -265
rect -1135 -271 -1131 -265
rect -1043 -266 -777 -265
rect -1425 -296 -1412 -271
rect -1381 -296 -1368 -271
rect -1212 -296 -1199 -271
rect -1168 -296 -1155 -271
rect -1486 -307 -1479 -303
rect -1459 -304 -1455 -296
rect -1459 -307 -1419 -304
rect -1469 -315 -1466 -311
rect -1459 -318 -1455 -307
rect -1447 -315 -1443 -310
rect -1423 -315 -1419 -307
rect -1415 -310 -1412 -296
rect -1371 -305 -1368 -296
rect -1371 -310 -1347 -305
rect -1340 -306 -1336 -296
rect -1415 -315 -1399 -310
rect -1379 -315 -1375 -311
rect -1415 -318 -1412 -315
rect -1371 -318 -1368 -310
rect -1340 -311 -1327 -306
rect -1340 -318 -1336 -311
rect -1273 -307 -1266 -303
rect -1246 -304 -1242 -296
rect -1246 -307 -1206 -304
rect -1256 -315 -1253 -311
rect -1246 -318 -1242 -307
rect -1234 -315 -1230 -310
rect -1210 -315 -1206 -307
rect -1202 -310 -1199 -296
rect -1158 -305 -1155 -296
rect -1158 -310 -1134 -305
rect -1127 -306 -1123 -296
rect -1015 -302 -1011 -266
rect -1202 -315 -1186 -310
rect -1166 -315 -1162 -311
rect -1202 -318 -1199 -315
rect -1158 -318 -1155 -310
rect -1127 -311 -1114 -306
rect -1127 -318 -1123 -311
rect -1467 -328 -1455 -318
rect -1423 -328 -1412 -318
rect -1379 -328 -1368 -318
rect -1254 -328 -1242 -318
rect -1210 -328 -1199 -318
rect -1166 -328 -1155 -318
rect -1479 -333 -1475 -328
rect -1443 -333 -1439 -328
rect -1399 -333 -1395 -328
rect -1348 -333 -1344 -328
rect -1266 -333 -1262 -328
rect -1230 -333 -1226 -328
rect -1186 -333 -1182 -328
rect -1135 -333 -1131 -328
rect -1480 -337 -1123 -333
rect -1127 -422 -1123 -337
rect -990 -334 -985 -279
rect -974 -298 -970 -291
rect -941 -298 -937 -291
rect -902 -303 -898 -266
rect -815 -286 -809 -279
rect -782 -282 -777 -266
rect -782 -283 -732 -282
rect -782 -285 -711 -283
rect -882 -291 -801 -286
rect -978 -334 -974 -330
rect -990 -338 -974 -334
rect -1024 -359 -1014 -354
rect -1007 -355 -1003 -342
rect -978 -350 -974 -338
rect -1007 -360 -994 -355
rect -1007 -362 -1003 -360
rect -970 -335 -966 -330
rect -970 -339 -953 -335
rect -970 -350 -966 -339
rect -957 -349 -953 -339
rect -945 -349 -941 -337
rect -957 -354 -941 -349
rect -1015 -421 -1011 -382
rect -974 -402 -970 -389
rect -957 -415 -951 -354
rect -945 -357 -941 -354
rect -937 -350 -933 -337
rect -937 -354 -916 -350
rect -937 -357 -933 -354
rect -922 -355 -916 -354
rect -922 -360 -912 -355
rect -906 -360 -901 -355
rect -894 -356 -890 -343
rect -852 -317 -843 -304
rect -804 -311 -801 -291
rect -769 -291 -766 -285
rect -750 -291 -747 -285
rect -735 -286 -711 -285
rect -729 -292 -726 -286
rect -760 -306 -757 -303
rect -760 -309 -747 -306
rect -804 -314 -768 -311
rect -750 -312 -747 -309
rect -750 -315 -728 -312
rect -720 -312 -717 -304
rect -365 -300 -361 150
rect -276 -149 -272 150
rect -213 -9 -209 150
rect -158 121 -154 150
rect 254 161 258 197
rect -115 139 -111 149
rect -77 139 -73 149
rect -33 139 -29 149
rect 5 139 9 149
rect -115 135 17 139
rect 279 129 284 184
rect 295 165 299 172
rect 328 165 332 172
rect 367 160 371 197
rect 414 177 465 183
rect 590 180 743 184
rect 387 172 465 177
rect 596 174 600 180
rect 634 174 638 180
rect 678 174 682 180
rect 723 174 727 180
rect 291 129 295 133
rect 279 125 295 129
rect -158 116 -53 121
rect -158 111 -154 116
rect -150 -9 -146 11
rect -80 110 -76 116
rect 245 104 255 109
rect 262 108 266 121
rect 291 113 295 125
rect 262 103 275 108
rect 262 101 266 103
rect 299 128 303 133
rect 299 124 316 128
rect 299 113 303 124
rect 312 114 316 124
rect 324 114 328 126
rect 312 109 328 114
rect 254 42 258 81
rect 295 61 299 74
rect 312 51 318 109
rect 324 106 328 109
rect 332 113 336 126
rect 646 149 659 174
rect 690 149 703 174
rect 575 138 592 142
rect 612 141 616 149
rect 612 138 652 141
rect 602 130 605 134
rect 612 127 616 138
rect 624 130 628 135
rect 648 130 652 138
rect 656 135 659 149
rect 700 140 703 149
rect 700 135 724 140
rect 731 139 735 149
rect 656 130 672 135
rect 692 130 696 134
rect 656 127 659 130
rect 700 127 703 135
rect 731 134 744 139
rect 731 127 735 134
rect 332 109 353 113
rect 332 106 336 109
rect 347 108 353 109
rect 347 103 357 108
rect 363 103 368 108
rect 375 107 379 120
rect 604 117 616 127
rect 648 117 659 127
rect 692 117 703 127
rect 592 112 596 117
rect 628 112 632 117
rect 672 112 676 117
rect 723 112 727 117
rect 591 108 735 112
rect 375 102 392 107
rect 375 100 379 102
rect 417 99 435 105
rect 328 61 332 74
rect 367 42 371 80
rect 417 62 425 99
rect 226 34 435 42
rect -213 -13 -142 -9
rect -213 -27 -209 -13
rect -205 -149 -201 -127
rect -150 -28 -146 -13
rect -276 -154 -197 -149
rect -276 -172 -272 -154
rect -205 -172 -201 -154
rect -268 -300 -264 -272
rect -365 -305 -259 -300
rect -720 -315 -708 -312
rect -852 -320 -758 -317
rect -894 -361 -877 -356
rect -894 -363 -890 -361
rect -941 -402 -937 -389
rect -902 -421 -898 -383
rect -852 -401 -844 -320
rect -750 -323 -747 -315
rect -720 -318 -717 -315
rect -365 -320 -361 -305
rect -268 -320 -264 -305
rect -729 -328 -726 -324
rect -739 -331 -711 -328
rect -769 -341 -766 -335
rect -739 -341 -735 -331
rect -834 -344 -735 -341
rect -834 -421 -823 -344
rect -1043 -422 -823 -421
rect -1127 -429 -823 -422
rect -357 -465 -353 -420
rect -1452 -575 -748 -571
rect -1446 -581 -1442 -575
rect -1408 -581 -1404 -575
rect -1364 -581 -1360 -575
rect -1319 -581 -1315 -575
rect -1233 -581 -1229 -575
rect -1195 -581 -1191 -575
rect -1151 -581 -1147 -575
rect -1106 -581 -1102 -575
rect -1014 -576 -748 -575
rect -1396 -606 -1383 -581
rect -1352 -606 -1339 -581
rect -1183 -606 -1170 -581
rect -1139 -606 -1126 -581
rect -1457 -617 -1450 -613
rect -1430 -614 -1426 -606
rect -1430 -617 -1390 -614
rect -1440 -625 -1437 -621
rect -1430 -628 -1426 -617
rect -1418 -625 -1414 -620
rect -1394 -625 -1390 -617
rect -1386 -620 -1383 -606
rect -1342 -615 -1339 -606
rect -1342 -620 -1318 -615
rect -1311 -616 -1307 -606
rect -1386 -625 -1370 -620
rect -1350 -625 -1346 -621
rect -1386 -628 -1383 -625
rect -1342 -628 -1339 -620
rect -1311 -621 -1298 -616
rect -1311 -628 -1307 -621
rect -1244 -617 -1237 -613
rect -1217 -614 -1213 -606
rect -1217 -617 -1177 -614
rect -1227 -625 -1224 -621
rect -1217 -628 -1213 -617
rect -1205 -625 -1201 -620
rect -1181 -625 -1177 -617
rect -1173 -620 -1170 -606
rect -1129 -615 -1126 -606
rect -1129 -620 -1105 -615
rect -1098 -616 -1094 -606
rect -986 -612 -982 -576
rect -1173 -625 -1157 -620
rect -1137 -625 -1133 -621
rect -1173 -628 -1170 -625
rect -1129 -628 -1126 -620
rect -1098 -621 -1085 -616
rect -1098 -628 -1094 -621
rect -1438 -638 -1426 -628
rect -1394 -638 -1383 -628
rect -1350 -638 -1339 -628
rect -1225 -638 -1213 -628
rect -1181 -638 -1170 -628
rect -1137 -638 -1126 -628
rect -1450 -643 -1446 -638
rect -1414 -643 -1410 -638
rect -1370 -643 -1366 -638
rect -1319 -643 -1315 -638
rect -1237 -643 -1233 -638
rect -1201 -643 -1197 -638
rect -1157 -643 -1153 -638
rect -1106 -643 -1102 -638
rect -1451 -647 -1094 -643
rect -1098 -732 -1094 -647
rect -961 -644 -956 -589
rect -945 -608 -941 -601
rect -912 -608 -908 -601
rect -873 -613 -869 -576
rect -786 -596 -780 -589
rect -753 -592 -748 -576
rect -349 -585 -345 -565
rect -260 -585 -256 -420
rect -197 -585 -193 -272
rect -142 -585 -138 -128
rect -72 -585 -68 10
rect 216 -111 449 -106
rect 244 -147 248 -111
rect 269 -179 274 -124
rect 285 -143 289 -136
rect 318 -143 322 -136
rect 357 -148 361 -111
rect 404 -131 455 -125
rect 580 -128 733 -124
rect 377 -136 455 -131
rect 586 -134 590 -128
rect 624 -134 628 -128
rect 668 -134 672 -128
rect 713 -134 717 -128
rect 281 -179 285 -175
rect 269 -183 285 -179
rect 235 -204 245 -199
rect 252 -200 256 -187
rect 281 -195 285 -183
rect 252 -205 265 -200
rect 252 -207 256 -205
rect 289 -180 293 -175
rect 289 -184 306 -180
rect 289 -195 293 -184
rect 302 -194 306 -184
rect 314 -194 318 -182
rect 302 -199 318 -194
rect 244 -266 248 -227
rect 285 -247 289 -234
rect 302 -257 308 -199
rect 314 -202 318 -199
rect 322 -195 326 -182
rect 636 -159 649 -134
rect 680 -159 693 -134
rect 565 -170 582 -166
rect 602 -167 606 -159
rect 602 -170 642 -167
rect 592 -178 595 -174
rect 602 -181 606 -170
rect 614 -178 618 -173
rect 638 -178 642 -170
rect 646 -173 649 -159
rect 690 -168 693 -159
rect 690 -173 714 -168
rect 721 -169 725 -159
rect 646 -178 662 -173
rect 682 -178 686 -174
rect 646 -181 649 -178
rect 690 -181 693 -173
rect 721 -174 734 -169
rect 721 -181 725 -174
rect 322 -199 343 -195
rect 322 -202 326 -199
rect 337 -200 343 -199
rect 337 -205 347 -200
rect 353 -205 358 -200
rect 365 -201 369 -188
rect 594 -191 606 -181
rect 638 -191 649 -181
rect 682 -191 693 -181
rect 582 -196 586 -191
rect 618 -196 622 -191
rect 662 -196 666 -191
rect 713 -196 717 -191
rect 581 -200 725 -196
rect 365 -206 382 -201
rect 365 -208 369 -206
rect 407 -209 425 -203
rect 318 -247 322 -234
rect 357 -266 361 -228
rect 407 -246 415 -209
rect 216 -274 425 -266
rect 240 -370 473 -365
rect 268 -406 272 -370
rect 293 -438 298 -383
rect 309 -402 313 -395
rect 342 -402 346 -395
rect 381 -407 385 -370
rect 428 -390 479 -384
rect 604 -387 757 -383
rect 401 -395 479 -390
rect 610 -393 614 -387
rect 648 -393 652 -387
rect 692 -393 696 -387
rect 737 -393 741 -387
rect 305 -438 309 -434
rect 293 -442 309 -438
rect 259 -463 269 -458
rect 276 -459 280 -446
rect 305 -454 309 -442
rect 276 -464 289 -459
rect 276 -466 280 -464
rect 313 -439 317 -434
rect 313 -443 330 -439
rect 313 -454 317 -443
rect 326 -453 330 -443
rect 338 -453 342 -441
rect 326 -458 342 -453
rect 268 -525 272 -486
rect 309 -506 313 -493
rect 326 -516 332 -458
rect 338 -461 342 -458
rect 346 -454 350 -441
rect 660 -418 673 -393
rect 704 -418 717 -393
rect 589 -429 606 -425
rect 626 -426 630 -418
rect 626 -429 666 -426
rect 616 -437 619 -433
rect 626 -440 630 -429
rect 638 -437 642 -432
rect 662 -437 666 -429
rect 670 -432 673 -418
rect 714 -427 717 -418
rect 714 -432 738 -427
rect 745 -428 749 -418
rect 670 -437 686 -432
rect 706 -437 710 -433
rect 670 -440 673 -437
rect 714 -440 717 -432
rect 745 -433 758 -428
rect 745 -440 749 -433
rect 346 -458 367 -454
rect 346 -461 350 -458
rect 361 -459 367 -458
rect 361 -464 371 -459
rect 377 -464 382 -459
rect 389 -460 393 -447
rect 618 -450 630 -440
rect 662 -450 673 -440
rect 706 -450 717 -440
rect 606 -455 610 -450
rect 642 -455 646 -450
rect 686 -455 690 -450
rect 737 -455 741 -450
rect 605 -459 749 -455
rect 389 -465 406 -460
rect 389 -467 393 -465
rect 431 -468 449 -462
rect 342 -506 346 -493
rect 381 -525 385 -487
rect 431 -505 439 -468
rect 240 -533 449 -525
rect -349 -589 -57 -585
rect -753 -593 -703 -592
rect -753 -595 -682 -593
rect -853 -601 -772 -596
rect -949 -644 -945 -640
rect -961 -648 -945 -644
rect -995 -669 -985 -664
rect -978 -665 -974 -652
rect -949 -660 -945 -648
rect -978 -670 -965 -665
rect -978 -672 -974 -670
rect -941 -645 -937 -640
rect -941 -649 -924 -645
rect -941 -660 -937 -649
rect -928 -659 -924 -649
rect -916 -659 -912 -647
rect -928 -664 -912 -659
rect -986 -731 -982 -692
rect -945 -712 -941 -699
rect -928 -725 -922 -664
rect -916 -667 -912 -664
rect -908 -660 -904 -647
rect -908 -664 -887 -660
rect -908 -667 -904 -664
rect -893 -665 -887 -664
rect -893 -670 -883 -665
rect -877 -670 -872 -665
rect -865 -666 -861 -653
rect -823 -627 -814 -614
rect -775 -621 -772 -601
rect -740 -601 -737 -595
rect -721 -601 -718 -595
rect -706 -596 -682 -595
rect -700 -602 -697 -596
rect -349 -598 -345 -589
rect -731 -616 -728 -613
rect -731 -619 -718 -616
rect -775 -624 -739 -621
rect -721 -622 -718 -619
rect -721 -625 -699 -622
rect -691 -622 -688 -614
rect -691 -625 -679 -622
rect -823 -630 -729 -627
rect -865 -671 -848 -666
rect -865 -673 -861 -671
rect -912 -712 -908 -699
rect -873 -731 -869 -693
rect -823 -711 -815 -630
rect -721 -633 -718 -625
rect -691 -628 -688 -625
rect -700 -638 -697 -634
rect -710 -641 -682 -638
rect -740 -651 -737 -645
rect -710 -651 -706 -641
rect -805 -654 -706 -651
rect -805 -731 -794 -654
rect 261 -676 494 -671
rect -341 -716 -337 -698
rect 289 -712 293 -676
rect -1014 -732 -794 -731
rect -1098 -739 -794 -732
rect 314 -744 319 -689
rect 330 -708 334 -701
rect 363 -708 367 -701
rect 402 -713 406 -676
rect 449 -696 500 -690
rect 625 -693 778 -689
rect 422 -701 500 -696
rect 631 -699 635 -693
rect 669 -699 673 -693
rect 713 -699 717 -693
rect 758 -699 762 -693
rect 326 -744 330 -740
rect 314 -748 330 -744
rect 280 -769 290 -764
rect 297 -765 301 -752
rect 326 -760 330 -748
rect 297 -770 310 -765
rect 297 -772 301 -770
rect 334 -745 338 -740
rect 334 -749 351 -745
rect 334 -760 338 -749
rect 347 -759 351 -749
rect 359 -759 363 -747
rect 347 -764 363 -759
rect 289 -831 293 -792
rect 330 -812 334 -799
rect 347 -822 353 -764
rect 359 -767 363 -764
rect 367 -760 371 -747
rect 681 -724 694 -699
rect 725 -724 738 -699
rect 610 -735 627 -731
rect 647 -732 651 -724
rect 647 -735 687 -732
rect 637 -743 640 -739
rect 647 -746 651 -735
rect 659 -743 663 -738
rect 683 -743 687 -735
rect 691 -738 694 -724
rect 735 -733 738 -724
rect 735 -738 759 -733
rect 766 -734 770 -724
rect 691 -743 707 -738
rect 727 -743 731 -739
rect 691 -746 694 -743
rect 735 -746 738 -738
rect 766 -739 779 -734
rect 766 -746 770 -739
rect 367 -764 388 -760
rect 367 -767 371 -764
rect 382 -765 388 -764
rect 382 -770 392 -765
rect 398 -770 403 -765
rect 410 -766 414 -753
rect 639 -756 651 -746
rect 683 -756 694 -746
rect 727 -756 738 -746
rect 627 -761 631 -756
rect 663 -761 667 -756
rect 707 -761 711 -756
rect 758 -761 762 -756
rect 626 -765 770 -761
rect 410 -771 427 -766
rect 410 -773 414 -771
rect 452 -774 470 -768
rect 363 -812 367 -799
rect 402 -831 406 -793
rect 452 -811 460 -774
rect 261 -839 470 -831
rect 690 -933 843 -929
rect 696 -939 700 -933
rect 734 -939 738 -933
rect 778 -939 782 -933
rect 823 -939 827 -933
rect 746 -964 759 -939
rect 790 -964 803 -939
rect 685 -975 692 -971
rect 712 -972 716 -964
rect 712 -975 752 -972
rect 702 -983 705 -979
rect 712 -986 716 -975
rect 724 -983 728 -978
rect 748 -983 752 -975
rect 756 -978 759 -964
rect 800 -973 803 -964
rect 800 -978 824 -973
rect 831 -974 835 -964
rect 756 -983 772 -978
rect 792 -983 796 -979
rect 756 -986 759 -983
rect 800 -986 803 -978
rect 831 -979 844 -974
rect 831 -986 835 -979
rect 704 -996 716 -986
rect 748 -996 759 -986
rect 792 -996 803 -986
rect 692 -1001 696 -996
rect 728 -1001 732 -996
rect 772 -1001 776 -996
rect 823 -1001 827 -996
rect 691 -1005 835 -1001
<< m2contact >>
rect -1366 284 -1355 291
rect -1029 317 -1023 322
rect -1153 284 -1142 291
rect -1013 305 -1008 310
rect -981 305 -976 310
rect -857 317 -847 324
rect -929 305 -921 310
rect -1068 237 -1063 242
rect -1033 236 -1027 241
rect -1013 189 -1008 194
rect -892 292 -881 298
rect -951 236 -945 241
rect -916 235 -910 240
rect -980 189 -975 194
rect -891 189 -883 195
rect -1351 -45 -1340 -38
rect -1014 -12 -1008 -7
rect -1138 -45 -1127 -38
rect -998 -24 -993 -19
rect -966 -24 -961 -19
rect -842 -12 -832 -5
rect -914 -24 -906 -19
rect -1053 -92 -1048 -87
rect -1018 -93 -1012 -88
rect -998 -140 -993 -135
rect -877 -37 -866 -31
rect -936 -93 -930 -88
rect -901 -94 -895 -89
rect -965 -140 -960 -135
rect -876 -140 -868 -134
rect -1327 -312 -1316 -305
rect -990 -279 -984 -274
rect -1114 -312 -1103 -305
rect -974 -291 -969 -286
rect -942 -291 -937 -286
rect -818 -279 -808 -272
rect -890 -291 -882 -286
rect -1029 -359 -1024 -354
rect -994 -360 -988 -355
rect -974 -407 -969 -402
rect -853 -304 -842 -298
rect -912 -360 -906 -355
rect 279 184 285 189
rect 295 172 300 177
rect 327 172 332 177
rect 379 172 387 177
rect 240 104 245 109
rect 275 103 281 108
rect 295 56 300 61
rect 570 137 575 142
rect 357 103 363 108
rect 392 102 398 107
rect 328 56 333 61
rect 312 45 318 51
rect 417 56 425 62
rect -877 -361 -871 -356
rect -941 -407 -936 -402
rect -852 -407 -844 -401
rect -1298 -622 -1287 -615
rect -961 -589 -955 -584
rect -1085 -622 -1074 -615
rect -945 -601 -940 -596
rect -913 -601 -908 -596
rect -789 -589 -779 -582
rect 269 -124 275 -119
rect 285 -136 290 -131
rect 317 -136 322 -131
rect 369 -136 377 -131
rect 230 -204 235 -199
rect 265 -205 271 -200
rect 285 -252 290 -247
rect 560 -171 565 -166
rect 347 -205 353 -200
rect 382 -206 388 -201
rect 318 -252 323 -247
rect 302 -263 308 -257
rect 407 -252 415 -246
rect 293 -383 299 -378
rect 309 -395 314 -390
rect 341 -395 346 -390
rect 393 -395 401 -390
rect 254 -463 259 -458
rect 289 -464 295 -459
rect 309 -511 314 -506
rect 584 -430 589 -425
rect 371 -464 377 -459
rect 406 -465 412 -460
rect 342 -511 347 -506
rect 326 -522 332 -516
rect 431 -511 439 -505
rect -861 -601 -853 -596
rect -1000 -669 -995 -664
rect -965 -670 -959 -665
rect -945 -717 -940 -712
rect -824 -614 -813 -608
rect -883 -670 -877 -665
rect -848 -671 -842 -666
rect -912 -717 -907 -712
rect -823 -717 -815 -711
rect 314 -689 320 -684
rect 330 -701 335 -696
rect 362 -701 367 -696
rect 414 -701 422 -696
rect 275 -769 280 -764
rect 310 -770 316 -765
rect 330 -817 335 -812
rect 605 -736 610 -731
rect 392 -770 398 -765
rect 427 -771 433 -766
rect 363 -817 368 -812
rect 347 -828 353 -822
rect 452 -817 460 -811
<< pm12contact >>
rect -115 172 -110 177
rect -77 172 -72 177
rect -33 172 -28 177
rect 5 172 10 177
rect -373 133 -368 138
rect -284 133 -279 138
rect -221 133 -216 138
rect -166 133 -161 138
rect -158 -1 -153 4
rect -80 -2 -75 3
rect -213 -139 -208 -134
rect -150 -140 -145 -135
rect -276 -284 -271 -279
rect -205 -284 -200 -279
rect -365 -432 -360 -427
rect -268 -432 -263 -427
rect -357 -577 -352 -572
rect -349 -710 -344 -705
<< metal2 >>
rect -1127 353 -1123 354
rect -1127 349 -849 353
rect -1340 338 -1145 342
rect -1340 290 -1336 338
rect -1355 285 -1336 290
rect -1127 290 -1123 349
rect -1084 340 -884 344
rect -1023 317 -910 322
rect -1142 285 -1123 290
rect -1068 305 -1013 310
rect -1008 305 -981 310
rect -976 305 -929 310
rect -1068 242 -1064 305
rect -1033 194 -1027 236
rect -951 195 -945 236
rect -916 240 -910 317
rect -890 298 -884 340
rect -854 324 -849 349
rect -1034 189 -1013 194
rect -1008 189 -980 194
rect -975 189 -961 194
rect -951 189 -891 195
rect 285 184 398 189
rect -118 172 -115 177
rect -80 172 -77 177
rect -36 172 -33 177
rect 2 172 5 177
rect 240 172 295 177
rect 300 172 327 177
rect 332 172 379 177
rect -377 133 -373 138
rect -288 133 -284 138
rect -225 133 -221 138
rect -170 133 -166 138
rect 240 109 244 172
rect 275 61 281 103
rect 357 62 363 103
rect 392 107 398 184
rect 274 56 295 61
rect 300 56 328 61
rect 333 56 347 61
rect 357 56 417 62
rect 570 49 575 137
rect 318 45 575 49
rect -1112 24 -1108 25
rect -1112 20 -834 24
rect -1325 9 -1130 13
rect -1325 -39 -1321 9
rect -1340 -44 -1321 -39
rect -1112 -39 -1108 20
rect -1069 11 -869 15
rect -1008 -12 -895 -7
rect -1127 -44 -1108 -39
rect -1053 -24 -998 -19
rect -993 -24 -966 -19
rect -961 -24 -914 -19
rect -1053 -87 -1049 -24
rect -1018 -135 -1012 -93
rect -936 -134 -930 -93
rect -901 -89 -895 -12
rect -875 -31 -869 11
rect -839 -5 -834 20
rect -163 -1 -158 4
rect -85 -2 -80 3
rect 275 -124 388 -119
rect -1019 -140 -998 -135
rect -993 -140 -965 -135
rect -960 -140 -946 -135
rect -936 -140 -876 -134
rect -218 -139 -213 -134
rect -155 -140 -150 -135
rect 230 -136 285 -131
rect 290 -136 317 -131
rect 322 -136 369 -131
rect 230 -199 234 -136
rect -1088 -243 -1084 -242
rect -1088 -247 -810 -243
rect 265 -247 271 -205
rect 347 -246 353 -205
rect 382 -201 388 -124
rect -1301 -258 -1106 -254
rect -1301 -306 -1297 -258
rect -1316 -311 -1297 -306
rect -1088 -306 -1084 -247
rect -1045 -256 -845 -252
rect -984 -279 -871 -274
rect -1103 -311 -1084 -306
rect -1029 -291 -974 -286
rect -969 -291 -942 -286
rect -937 -291 -890 -286
rect -1029 -354 -1025 -291
rect -994 -402 -988 -360
rect -912 -401 -906 -360
rect -877 -356 -871 -279
rect -851 -298 -845 -256
rect -815 -272 -810 -247
rect 264 -252 285 -247
rect 290 -252 318 -247
rect 323 -252 337 -247
rect 347 -252 407 -246
rect 560 -259 565 -171
rect 308 -263 565 -259
rect -281 -284 -276 -279
rect -210 -284 -205 -279
rect 299 -383 412 -378
rect 254 -395 309 -390
rect 314 -395 341 -390
rect 346 -395 393 -390
rect -995 -407 -974 -402
rect -969 -407 -941 -402
rect -936 -407 -922 -402
rect -912 -407 -852 -401
rect -370 -432 -365 -427
rect -273 -432 -268 -427
rect 254 -458 258 -395
rect 289 -506 295 -464
rect 371 -505 377 -464
rect 406 -460 412 -383
rect 288 -511 309 -506
rect 314 -511 342 -506
rect 347 -511 361 -506
rect 371 -511 431 -505
rect 584 -518 589 -430
rect 332 -522 589 -518
rect -1059 -553 -1055 -552
rect -1059 -557 -781 -553
rect -1272 -568 -1077 -564
rect -1272 -616 -1268 -568
rect -1287 -621 -1268 -616
rect -1059 -616 -1055 -557
rect -1016 -566 -816 -562
rect -955 -589 -842 -584
rect -1074 -621 -1055 -616
rect -1000 -601 -945 -596
rect -940 -601 -913 -596
rect -908 -601 -861 -596
rect -1000 -664 -996 -601
rect -965 -712 -959 -670
rect -883 -711 -877 -670
rect -848 -666 -842 -589
rect -822 -608 -816 -566
rect -786 -582 -781 -557
rect -362 -577 -357 -572
rect 320 -689 433 -684
rect 275 -701 330 -696
rect 335 -701 362 -696
rect 367 -701 414 -696
rect -354 -710 -349 -705
rect -966 -717 -945 -712
rect -940 -717 -912 -712
rect -907 -717 -893 -712
rect -883 -717 -823 -711
rect 275 -764 279 -701
rect 310 -812 316 -770
rect 392 -811 398 -770
rect 427 -766 433 -689
rect 309 -817 330 -812
rect 335 -817 363 -812
rect 368 -817 382 -812
rect 392 -817 452 -811
rect 605 -824 610 -736
rect 353 -828 610 -824
<< m3contact >>
rect -1145 337 -1132 343
rect -1094 338 -1084 344
rect -1130 8 -1117 14
rect -1079 9 -1069 15
rect -1106 -259 -1093 -253
rect -1055 -258 -1045 -252
rect -1077 -569 -1064 -563
rect -1026 -568 -1016 -562
<< metal3 >>
rect -1132 338 -1094 343
rect -1117 9 -1079 14
rect -1093 -258 -1055 -253
rect -1064 -568 -1026 -563
<< labels >>
rlabel metal1 -166 215 -162 219 5 vdd!
rlabel metal2 -170 133 -167 138 1 u1
rlabel metal1 -146 -13 -142 -9 1 r3
rlabel metal1 -221 215 -217 219 5 vdd!
rlabel metal2 -225 133 -222 138 1 u1
rlabel metal1 -201 -154 -197 -149 1 r2
rlabel metal1 -284 215 -280 219 5 vdd!
rlabel metal2 -288 133 -285 138 1 u1
rlabel metal1 -76 116 -53 121 1 r4
rlabel metal1 -264 -305 -259 -300 1 r1
rlabel metal1 -373 215 -369 219 5 vdd!
rlabel metal2 -377 133 -374 138 2 u1
rlabel metal1 -365 137 -361 141 1 r1
rlabel metal1 -341 -716 -337 -712 1 gnd!
rlabel metal2 -354 -710 -350 -705 1 u1
rlabel metal1 -121 240 23 245 5 vdd!
rlabel metal1 -115 135 17 139 1 gnd!
rlabel metal2 -118 172 -115 177 1 r1
rlabel metal2 -80 172 -77 177 1 r2
rlabel metal2 -36 172 -33 177 1 r3
rlabel metal2 2 172 5 177 1 r4
rlabel metal1 -107 172 -103 177 1 c0
rlabel metal1 -69 171 -65 177 1 c1
rlabel metal1 -25 171 -21 177 1 c2
rlabel metal1 13 171 17 177 1 out_carry
rlabel metal2 -362 -577 -358 -572 1 carry_reg
rlabel metal2 -370 -432 -366 -427 1 p0
rlabel metal2 -273 -432 -269 -427 1 g0
rlabel metal2 -281 -284 -277 -279 1 p1
rlabel metal2 -210 -284 -206 -279 1 g1
rlabel metal2 -218 -139 -214 -134 1 p2
rlabel metal2 -155 -140 -151 -135 1 g2
rlabel metal2 -163 -1 -159 4 1 p3
rlabel metal2 -85 -2 -81 3 1 g3
rlabel metal1 -752 281 -747 284 1 g0
rlabel metal1 -814 276 -811 279 1 b0_reg
rlabel metal1 -814 282 -810 285 1 a0_reg
rlabel metal1 -996 182 -990 188 1 p0
rlabel metal1 -997 168 -883 174 1 gnd
rlabel metal1 -1295 282 -1293 284 1 clk
rlabel metal1 -1297 261 -1294 262 1 gnd
rlabel metal1 -1291 333 -1289 334 5 vdd
rlabel metal1 -1272 282 -1271 284 1 clk
rlabel metal1 -1204 282 -1202 284 1 clk
rlabel metal1 -1160 287 -1157 289 1 a0_reg
rlabel metal1 -1310 290 -1308 292 3 a0
rlabel metal1 -1417 282 -1415 284 1 clk
rlabel metal1 -1485 282 -1484 284 1 clk
rlabel metal1 -1504 333 -1502 334 5 vdd
rlabel metal1 -1510 261 -1507 262 1 gnd
rlabel metal1 -1508 282 -1506 284 1 clk
rlabel metal1 -1523 290 -1521 292 3 b0
rlabel metal1 -1373 287 -1370 289 1 b0_reg
rlabel metal1 -982 -161 -868 -155 1 gnd
rlabel metal1 -1280 -47 -1278 -45 1 clk
rlabel metal1 -1282 -68 -1279 -67 1 gnd
rlabel metal1 -1276 4 -1274 5 5 vdd
rlabel metal1 -1257 -47 -1256 -45 1 clk
rlabel metal1 -1189 -47 -1187 -45 1 clk
rlabel metal1 -1402 -47 -1400 -45 1 clk
rlabel metal1 -1470 -47 -1469 -45 1 clk
rlabel metal1 -1489 4 -1487 5 5 vdd
rlabel metal1 -1495 -68 -1492 -67 1 gnd
rlabel metal1 -1493 -47 -1491 -45 1 clk
rlabel metal1 -958 -428 -844 -422 1 gnd
rlabel metal1 -1256 -314 -1254 -312 1 clk
rlabel metal1 -1258 -335 -1255 -334 1 gnd
rlabel metal1 -1252 -263 -1250 -262 5 vdd
rlabel metal1 -1233 -314 -1232 -312 1 clk
rlabel metal1 -1165 -314 -1163 -312 1 clk
rlabel metal1 -1378 -314 -1376 -312 1 clk
rlabel metal1 -1446 -314 -1445 -312 1 clk
rlabel metal1 -1465 -263 -1463 -262 5 vdd
rlabel metal1 -1471 -335 -1468 -334 1 gnd
rlabel metal1 -1469 -314 -1467 -312 1 clk
rlabel metal1 -1440 -624 -1438 -622 1 clk
rlabel metal1 -1442 -645 -1439 -644 1 gnd
rlabel metal1 -1436 -573 -1434 -572 5 vdd
rlabel metal1 -1417 -624 -1416 -622 1 clk
rlabel metal1 -1349 -624 -1347 -622 1 clk
rlabel metal1 -1136 -624 -1134 -622 1 clk
rlabel metal1 -1204 -624 -1203 -622 1 clk
rlabel metal1 -1223 -573 -1221 -572 5 vdd
rlabel metal1 -1229 -645 -1226 -644 1 gnd
rlabel metal1 -1227 -624 -1225 -622 1 clk
rlabel metal1 -929 -738 -815 -732 1 gnd
rlabel metal1 -1295 -39 -1293 -37 1 a1
rlabel metal1 -1360 -42 -1355 -40 1 b1_reg
rlabel metal1 -1508 -39 -1506 -37 1 b1
rlabel metal1 -1145 -42 -1142 -40 1 a1_reg
rlabel metal1 -981 -147 -975 -141 1 p1
rlabel metal1 -799 -53 -796 -50 1 b1_reg
rlabel metal1 -799 -47 -795 -44 1 a1_reg
rlabel metal1 -737 -48 -732 -45 1 g1
rlabel metal1 -1271 -306 -1269 -304 1 a2
rlabel metal1 -1121 -309 -1118 -307 1 a2_reg
rlabel metal1 -1334 -309 -1331 -307 1 b2_reg
rlabel metal1 -1484 -306 -1481 -304 1 b2
rlabel metal1 -775 -314 -771 -311 1 a2_reg
rlabel metal1 -775 -320 -771 -317 1 b2_reg
rlabel metal1 -957 -414 -951 -408 1 p2
rlabel metal1 -713 -315 -708 -312 1 g2
rlabel metal1 -684 -625 -679 -622 7 g3
rlabel metal1 -746 -624 -741 -621 1 a3_reg
rlabel metal1 -746 -630 -741 -627 1 b3_reg
rlabel metal1 -928 -724 -922 -718 1 p3
rlabel metal1 -1092 -619 -1089 -617 1 a3_reg
rlabel metal1 -1242 -616 -1239 -614 1 a3
rlabel metal1 -1305 -619 -1302 -617 1 b3_reg
rlabel metal1 -1455 -616 -1452 -614 1 b3
rlabel metal1 -583 -11 -583 -11 5 vdd!
rlabel metal1 -577 -56 -577 -56 1 gnd!
rlabel metal1 -597 -41 -594 -38 1 clk
rlabel metal1 -576 -41 -573 -38 1 u1
rlabel metal1 -634 252 -632 254 3 carry
rlabel metal1 -485 249 -480 251 1 carry_reg
rlabel metal1 -528 244 -526 246 1 clk
rlabel metal1 -596 244 -595 246 1 clk
rlabel metal1 -615 295 -613 296 5 vdd
rlabel metal1 -621 223 -618 224 1 gnd
rlabel metal1 -619 244 -617 246 1 clk
rlabel metal1 423 178 460 183 1 carry_reg
rlabel metal1 458 -695 495 -690 1 c2
rlabel metal1 452 -774 468 -768 1 p3
rlabel metal1 437 -389 474 -384 1 c1
rlabel metal1 431 -468 447 -462 1 p2
rlabel metal1 407 -209 423 -203 1 p1
rlabel metal1 413 -130 450 -125 1 c0
rlabel metal1 622 -734 624 -732 1 s3
rlabel metal1 772 -737 775 -735 1 s3_reg
rlabel metal1 751 -431 754 -429 1 s2_reg
rlabel metal1 601 -428 603 -426 1 s2
rlabel metal1 347 -821 353 -817 1 s3
rlabel metal1 326 -515 332 -511 1 s2
rlabel metal1 302 -256 308 -252 1 s1
rlabel metal1 727 -172 730 -170 1 s1_reg
rlabel metal1 577 -169 579 -167 1 s1
rlabel metal1 637 -742 639 -740 1 clk
rlabel metal1 635 -763 638 -762 1 gnd
rlabel metal1 641 -691 643 -690 5 vdd
rlabel metal1 660 -742 661 -740 1 clk
rlabel metal1 728 -742 730 -740 1 clk
rlabel metal1 370 -676 484 -671 5 VDD
rlabel metal1 346 -838 460 -832 1 GND
rlabel metal1 836 -977 841 -975 1 out_carry_reg
rlabel metal1 687 -974 689 -972 1 out_carry
rlabel metal1 793 -982 795 -980 1 clk
rlabel metal1 725 -982 726 -980 1 clk
rlabel metal1 706 -931 708 -930 5 vdd
rlabel metal1 700 -1003 703 -1002 1 gnd
rlabel metal1 702 -982 704 -980 1 clk
rlabel metal1 616 -436 618 -434 1 clk
rlabel metal1 614 -457 617 -456 1 gnd
rlabel metal1 620 -385 622 -384 5 vdd
rlabel metal1 639 -436 640 -434 1 clk
rlabel metal1 707 -436 709 -434 1 clk
rlabel metal1 349 -370 463 -365 5 VDD
rlabel metal1 325 -532 439 -526 1 GND
rlabel metal1 592 -177 594 -175 1 clk
rlabel metal1 590 -198 593 -197 1 gnd
rlabel metal1 596 -126 598 -125 5 vdd
rlabel metal1 615 -177 616 -175 1 clk
rlabel metal1 683 -177 685 -175 1 clk
rlabel metal1 325 -111 439 -106 5 VDD
rlabel metal1 301 -273 415 -267 1 GND
rlabel metal1 312 52 318 56 1 s0
rlabel metal1 587 139 589 141 1 s0
rlabel metal1 737 136 740 138 1 s0_reg
rlabel metal1 602 131 604 133 1 clk
rlabel metal1 600 110 603 111 1 gnd
rlabel metal1 606 182 608 183 5 vdd
rlabel metal1 625 131 626 133 1 clk
rlabel metal1 693 131 695 133 1 clk
rlabel metal1 417 99 433 105 1 p0
rlabel metal1 335 197 449 202 5 VDD
rlabel metal1 311 35 425 41 1 GND
<< end >>
