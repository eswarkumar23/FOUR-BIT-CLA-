magic
tech scmos
timestamp 1731668181
<< nwell >>
rect 0 0 34 36
rect 41 -1 65 23
<< polysilicon >>
rect 11 30 13 33
rect 21 30 23 33
rect 52 17 54 20
rect 11 -15 13 6
rect 21 -15 23 6
rect 52 -9 54 5
rect 52 -18 54 -15
rect 11 -24 13 -21
rect 21 -24 23 -21
<< ndiffusion >>
rect 51 -15 52 -9
rect 54 -15 55 -9
rect 10 -21 11 -15
rect 13 -21 15 -15
rect 19 -21 21 -15
rect 23 -21 24 -15
<< pdiffusion >>
rect 10 6 11 30
rect 13 6 21 30
rect 23 6 24 30
rect 51 5 52 17
rect 54 5 55 17
<< metal1 >>
rect 0 36 42 39
rect 6 30 9 36
rect 39 26 42 36
rect 39 23 65 26
rect 0 -5 17 -2
rect 25 -3 28 6
rect 47 17 50 23
rect 25 -6 48 -3
rect 56 -3 59 5
rect 56 -6 65 -3
rect 0 -11 7 -8
rect 25 -9 28 -6
rect 56 -9 59 -6
rect 16 -12 28 -9
rect 16 -15 19 -12
rect 47 -19 50 -15
rect 6 -27 9 -21
rect 25 -27 28 -21
rect 37 -22 65 -19
rect 37 -27 41 -22
rect 0 -30 41 -27
<< ntransistor >>
rect 52 -15 54 -9
rect 11 -21 13 -15
rect 21 -21 23 -15
<< ptransistor >>
rect 11 6 13 30
rect 21 6 23 30
rect 52 5 54 17
<< polycontact >>
rect 7 -12 11 -8
rect 17 -5 21 -1
rect 48 -6 52 -2
<< ndcontact >>
rect 47 -15 51 -9
rect 55 -15 59 -9
rect 6 -21 10 -15
rect 15 -21 19 -15
rect 24 -21 28 -15
<< pdcontact >>
rect 6 6 10 30
rect 24 6 28 30
rect 47 5 51 17
rect 55 5 59 17
<< labels >>
rlabel metal1 18 37 18 37 5 vdd!
rlabel metal1 34 -6 34 -3 7 out
rlabel metal1 21 -28 21 -28 1 gnd!
rlabel metal1 0 -5 0 -2 3 b
rlabel metal1 0 -11 0 -8 3 a
rlabel metal1 55 24 55 24 5 vdd!
rlabel metal1 61 -21 61 -21 1 gnd!
rlabel metal1 65 -6 65 -3 7 op
rlabel metal1 41 -6 41 -3 3 in
<< end >>
