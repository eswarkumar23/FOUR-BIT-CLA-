magic
tech scmos
timestamp 1732055747
<< nwell >>
rect 254 -29 279 28
rect 291 -57 316 -17
rect 324 -24 349 16
rect 367 -30 392 27
rect 500 14 534 38
rect 540 13 564 37
<< ntransistor >>
rect 302 -7 304 13
rect 511 -12 513 0
rect 521 -12 523 0
rect 551 -1 553 5
rect 265 -59 267 -39
rect 335 -54 337 -34
rect 378 -60 380 -40
<< ptransistor >>
rect 265 -19 267 21
rect 511 20 513 32
rect 521 20 523 32
rect 335 -14 337 6
rect 378 -20 380 20
rect 551 19 553 31
rect 302 -47 304 -27
<< ndiffusion >>
rect 301 -7 302 13
rect 304 -7 305 13
rect 510 -12 511 0
rect 513 -12 521 0
rect 523 -12 524 0
rect 550 -1 551 5
rect 553 -1 554 5
rect 264 -59 265 -39
rect 267 -59 268 -39
rect 334 -54 335 -34
rect 337 -54 338 -34
rect 377 -60 378 -40
rect 380 -60 381 -40
<< pdiffusion >>
rect 264 -19 265 21
rect 267 -19 268 21
rect 510 20 511 32
rect 513 20 515 32
rect 519 20 521 32
rect 523 20 524 32
rect 334 -14 335 6
rect 337 -14 338 6
rect 377 -20 378 20
rect 380 -20 381 20
rect 550 19 551 31
rect 553 19 554 31
rect 301 -47 302 -27
rect 304 -47 305 -27
<< ndcontact >>
rect 297 -7 301 13
rect 305 -7 309 13
rect 506 -12 510 0
rect 524 -12 528 0
rect 546 -1 550 5
rect 554 -1 558 5
rect 260 -59 264 -39
rect 268 -59 272 -39
rect 330 -54 334 -34
rect 338 -54 342 -34
rect 373 -60 377 -40
rect 381 -60 385 -40
<< pdcontact >>
rect 260 -19 264 21
rect 268 -19 272 21
rect 506 20 510 32
rect 515 20 519 32
rect 524 20 528 32
rect 330 -14 334 6
rect 338 -14 342 6
rect 373 -20 377 20
rect 381 -20 385 20
rect 546 19 550 31
rect 554 19 558 31
rect 297 -47 301 -27
rect 305 -47 309 -27
<< polysilicon >>
rect 511 32 513 35
rect 521 32 523 35
rect 265 21 267 25
rect 378 20 380 24
rect 551 31 553 34
rect 302 13 304 20
rect 335 6 337 20
rect 302 -10 304 -7
rect 335 -17 337 -14
rect 265 -39 267 -19
rect 511 0 513 20
rect 521 0 523 20
rect 551 5 553 19
rect 551 -4 553 -1
rect 511 -15 513 -12
rect 521 -15 523 -12
rect 302 -27 304 -24
rect 335 -34 337 -31
rect 265 -62 267 -59
rect 302 -61 304 -47
rect 378 -40 380 -20
rect 335 -61 337 -54
rect 378 -63 380 -60
<< polycontact >>
rect 301 20 305 25
rect 334 20 338 25
rect 261 -36 265 -31
rect 507 9 511 13
rect 517 3 521 7
rect 547 8 551 12
rect 374 -37 378 -32
rect 301 -66 305 -61
rect 334 -66 338 -61
<< metal1 >>
rect 232 57 498 62
rect 260 21 264 57
rect 285 -11 290 44
rect 301 25 305 32
rect 334 25 338 32
rect 373 20 377 57
rect 493 41 498 57
rect 493 40 543 41
rect 493 38 564 40
rect 393 32 474 37
rect 297 -11 301 -7
rect 285 -15 301 -11
rect 251 -36 261 -31
rect 268 -32 272 -19
rect 297 -27 301 -15
rect 268 -37 281 -32
rect 268 -39 272 -37
rect 305 -12 309 -7
rect 305 -16 322 -12
rect 305 -27 309 -16
rect 318 -26 322 -16
rect 330 -26 334 -14
rect 318 -31 334 -26
rect 260 -98 264 -59
rect 301 -79 305 -66
rect 318 -92 324 -31
rect 330 -34 334 -31
rect 338 -27 342 -14
rect 471 12 474 32
rect 506 32 509 38
rect 525 32 528 38
rect 540 37 564 38
rect 546 31 549 37
rect 515 17 518 20
rect 515 14 528 17
rect 471 9 507 12
rect 525 11 528 14
rect 525 8 547 11
rect 555 11 558 19
rect 555 8 567 11
rect 338 -31 359 -27
rect 338 -34 342 -31
rect 353 -32 359 -31
rect 353 -37 363 -32
rect 369 -37 374 -32
rect 381 -33 385 -20
rect 423 3 517 6
rect 381 -38 398 -33
rect 381 -40 385 -38
rect 334 -79 338 -66
rect 373 -98 377 -60
rect 423 -78 431 3
rect 525 0 528 8
rect 555 5 558 8
rect 546 -5 549 -1
rect 536 -8 564 -5
rect 506 -18 509 -12
rect 536 -18 540 -8
rect 441 -21 540 -18
rect 441 -98 452 -21
rect 232 -106 452 -98
<< m2contact >>
rect 285 44 291 49
rect 301 32 306 37
rect 333 32 338 37
rect 385 32 393 37
rect 246 -36 251 -31
rect 281 -37 287 -32
rect 301 -84 306 -79
rect 363 -37 369 -32
rect 398 -38 404 -33
rect 334 -84 339 -79
rect 423 -84 431 -78
<< metal2 >>
rect 291 44 404 49
rect 246 32 301 37
rect 306 32 333 37
rect 338 32 385 37
rect 246 -31 250 32
rect 281 -79 287 -37
rect 363 -78 369 -37
rect 398 -33 404 44
rect 280 -84 301 -79
rect 306 -84 334 -79
rect 339 -84 353 -79
rect 363 -84 423 -78
<< labels >>
rlabel metal1 562 8 567 11 1 g0
rlabel metal1 500 3 503 6 1 b0_reg
rlabel metal1 500 9 504 12 1 a0_reg
rlabel metal1 560 -7 560 -7 1 gnd!
rlabel metal1 554 38 554 38 5 vdd!
rlabel metal1 534 8 534 11 7 out
rlabel metal1 524 -20 524 -20 1 gnd!
rlabel metal1 524 40 524 40 5 vdd!
rlabel metal1 457 32 472 37 1 a0_reg
rlabel metal1 423 -19 431 -3 1 b0_reg
rlabel metal1 318 -91 324 -85 1 p0
rlabel metal1 341 57 455 62 1 vdd
rlabel metal1 317 -105 431 -99 1 gnd
<< end >>
