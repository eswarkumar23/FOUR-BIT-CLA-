magic
tech scmos
timestamp 1732056734
<< nwell >>
rect -392 -175 -360 -138
rect -354 -175 -328 -138
rect -310 -175 -284 -138
rect -265 -175 -239 -138
rect -113 -243 -88 -186
rect -76 -271 -51 -231
rect -43 -238 -18 -198
rect 0 -244 25 -187
rect 229 -211 261 -174
rect 267 -211 293 -174
rect 311 -211 337 -174
rect 356 -211 382 -174
rect -123 -551 -98 -494
rect -86 -579 -61 -539
rect -53 -546 -28 -506
rect -10 -552 15 -495
rect 219 -519 251 -482
rect 257 -519 283 -482
rect 301 -519 327 -482
rect 346 -519 372 -482
rect -99 -810 -74 -753
rect -62 -838 -37 -798
rect -29 -805 -4 -765
rect 14 -811 39 -754
rect 243 -778 275 -741
rect 281 -778 307 -741
rect 325 -778 351 -741
rect 370 -778 396 -741
rect -78 -1116 -53 -1059
rect -41 -1144 -16 -1104
rect -8 -1111 17 -1071
rect 35 -1117 60 -1060
rect 264 -1084 296 -1047
rect 302 -1084 328 -1047
rect 346 -1084 372 -1047
rect 391 -1084 417 -1047
rect 329 -1324 361 -1287
rect 367 -1324 393 -1287
rect 411 -1324 437 -1287
rect 456 -1324 482 -1287
<< ntransistor >>
rect -385 -201 -383 -191
rect -349 -201 -347 -191
rect -341 -201 -339 -191
rect -305 -201 -303 -191
rect -297 -201 -295 -191
rect -254 -201 -252 -191
rect -65 -221 -63 -201
rect -102 -273 -100 -253
rect -32 -268 -30 -248
rect 236 -237 238 -227
rect 272 -237 274 -227
rect 280 -237 282 -227
rect 316 -237 318 -227
rect 324 -237 326 -227
rect 367 -237 369 -227
rect 11 -274 13 -254
rect -75 -529 -73 -509
rect -112 -581 -110 -561
rect -42 -576 -40 -556
rect 226 -545 228 -535
rect 262 -545 264 -535
rect 270 -545 272 -535
rect 306 -545 308 -535
rect 314 -545 316 -535
rect 357 -545 359 -535
rect 1 -582 3 -562
rect -51 -788 -49 -768
rect -88 -840 -86 -820
rect -18 -835 -16 -815
rect 250 -804 252 -794
rect 286 -804 288 -794
rect 294 -804 296 -794
rect 330 -804 332 -794
rect 338 -804 340 -794
rect 381 -804 383 -794
rect 25 -841 27 -821
rect -30 -1094 -28 -1074
rect -67 -1146 -65 -1126
rect 3 -1141 5 -1121
rect 271 -1110 273 -1100
rect 307 -1110 309 -1100
rect 315 -1110 317 -1100
rect 351 -1110 353 -1100
rect 359 -1110 361 -1100
rect 402 -1110 404 -1100
rect 46 -1147 48 -1127
rect 336 -1350 338 -1340
rect 372 -1350 374 -1340
rect 380 -1350 382 -1340
rect 416 -1350 418 -1340
rect 424 -1350 426 -1340
rect 467 -1350 469 -1340
<< ptransistor >>
rect -381 -169 -379 -144
rect -373 -169 -371 -144
rect -343 -169 -341 -144
rect -299 -169 -297 -144
rect -254 -169 -252 -144
rect -102 -233 -100 -193
rect -32 -228 -30 -208
rect 11 -234 13 -194
rect 240 -205 242 -180
rect 248 -205 250 -180
rect 278 -205 280 -180
rect 322 -205 324 -180
rect 367 -205 369 -180
rect -65 -261 -63 -241
rect -112 -541 -110 -501
rect -42 -536 -40 -516
rect 1 -542 3 -502
rect 230 -513 232 -488
rect 238 -513 240 -488
rect 268 -513 270 -488
rect 312 -513 314 -488
rect 357 -513 359 -488
rect -75 -569 -73 -549
rect -88 -800 -86 -760
rect -18 -795 -16 -775
rect 25 -801 27 -761
rect 254 -772 256 -747
rect 262 -772 264 -747
rect 292 -772 294 -747
rect 336 -772 338 -747
rect 381 -772 383 -747
rect -51 -828 -49 -808
rect -67 -1106 -65 -1066
rect 3 -1101 5 -1081
rect 46 -1107 48 -1067
rect 275 -1078 277 -1053
rect 283 -1078 285 -1053
rect 313 -1078 315 -1053
rect 357 -1078 359 -1053
rect 402 -1078 404 -1053
rect -30 -1134 -28 -1114
rect 340 -1318 342 -1293
rect 348 -1318 350 -1293
rect 378 -1318 380 -1293
rect 422 -1318 424 -1293
rect 467 -1318 469 -1293
<< ndiffusion >>
rect -386 -201 -385 -191
rect -383 -201 -382 -191
rect -350 -201 -349 -191
rect -347 -201 -346 -191
rect -342 -201 -341 -191
rect -339 -201 -338 -191
rect -306 -201 -305 -191
rect -303 -201 -302 -191
rect -298 -201 -297 -191
rect -295 -201 -294 -191
rect -255 -201 -254 -191
rect -252 -201 -251 -191
rect -66 -221 -65 -201
rect -63 -221 -62 -201
rect -103 -273 -102 -253
rect -100 -273 -99 -253
rect -33 -268 -32 -248
rect -30 -268 -29 -248
rect 235 -237 236 -227
rect 238 -237 239 -227
rect 271 -237 272 -227
rect 274 -237 275 -227
rect 279 -237 280 -227
rect 282 -237 283 -227
rect 315 -237 316 -227
rect 318 -237 319 -227
rect 323 -237 324 -227
rect 326 -237 327 -227
rect 366 -237 367 -227
rect 369 -237 370 -227
rect 10 -274 11 -254
rect 13 -274 14 -254
rect -76 -529 -75 -509
rect -73 -529 -72 -509
rect -113 -581 -112 -561
rect -110 -581 -109 -561
rect -43 -576 -42 -556
rect -40 -576 -39 -556
rect 225 -545 226 -535
rect 228 -545 229 -535
rect 261 -545 262 -535
rect 264 -545 265 -535
rect 269 -545 270 -535
rect 272 -545 273 -535
rect 305 -545 306 -535
rect 308 -545 309 -535
rect 313 -545 314 -535
rect 316 -545 317 -535
rect 356 -545 357 -535
rect 359 -545 360 -535
rect 0 -582 1 -562
rect 3 -582 4 -562
rect -52 -788 -51 -768
rect -49 -788 -48 -768
rect -89 -840 -88 -820
rect -86 -840 -85 -820
rect -19 -835 -18 -815
rect -16 -835 -15 -815
rect 249 -804 250 -794
rect 252 -804 253 -794
rect 285 -804 286 -794
rect 288 -804 289 -794
rect 293 -804 294 -794
rect 296 -804 297 -794
rect 329 -804 330 -794
rect 332 -804 333 -794
rect 337 -804 338 -794
rect 340 -804 341 -794
rect 380 -804 381 -794
rect 383 -804 384 -794
rect 24 -841 25 -821
rect 27 -841 28 -821
rect -31 -1094 -30 -1074
rect -28 -1094 -27 -1074
rect -68 -1146 -67 -1126
rect -65 -1146 -64 -1126
rect 2 -1141 3 -1121
rect 5 -1141 6 -1121
rect 270 -1110 271 -1100
rect 273 -1110 274 -1100
rect 306 -1110 307 -1100
rect 309 -1110 310 -1100
rect 314 -1110 315 -1100
rect 317 -1110 318 -1100
rect 350 -1110 351 -1100
rect 353 -1110 354 -1100
rect 358 -1110 359 -1100
rect 361 -1110 362 -1100
rect 401 -1110 402 -1100
rect 404 -1110 405 -1100
rect 45 -1147 46 -1127
rect 48 -1147 49 -1127
rect 335 -1350 336 -1340
rect 338 -1350 339 -1340
rect 371 -1350 372 -1340
rect 374 -1350 375 -1340
rect 379 -1350 380 -1340
rect 382 -1350 383 -1340
rect 415 -1350 416 -1340
rect 418 -1350 419 -1340
rect 423 -1350 424 -1340
rect 426 -1350 427 -1340
rect 466 -1350 467 -1340
rect 469 -1350 470 -1340
<< pdiffusion >>
rect -382 -169 -381 -144
rect -379 -169 -378 -144
rect -374 -169 -373 -144
rect -371 -169 -370 -144
rect -344 -169 -343 -144
rect -341 -169 -340 -144
rect -300 -169 -299 -144
rect -297 -169 -296 -144
rect -255 -169 -254 -144
rect -252 -169 -251 -144
rect -103 -233 -102 -193
rect -100 -233 -99 -193
rect -33 -228 -32 -208
rect -30 -228 -29 -208
rect 10 -234 11 -194
rect 13 -234 14 -194
rect 239 -205 240 -180
rect 242 -205 243 -180
rect 247 -205 248 -180
rect 250 -205 251 -180
rect 277 -205 278 -180
rect 280 -205 281 -180
rect 321 -205 322 -180
rect 324 -205 325 -180
rect 366 -205 367 -180
rect 369 -205 370 -180
rect -66 -261 -65 -241
rect -63 -261 -62 -241
rect -113 -541 -112 -501
rect -110 -541 -109 -501
rect -43 -536 -42 -516
rect -40 -536 -39 -516
rect 0 -542 1 -502
rect 3 -542 4 -502
rect 229 -513 230 -488
rect 232 -513 233 -488
rect 237 -513 238 -488
rect 240 -513 241 -488
rect 267 -513 268 -488
rect 270 -513 271 -488
rect 311 -513 312 -488
rect 314 -513 315 -488
rect 356 -513 357 -488
rect 359 -513 360 -488
rect -76 -569 -75 -549
rect -73 -569 -72 -549
rect -89 -800 -88 -760
rect -86 -800 -85 -760
rect -19 -795 -18 -775
rect -16 -795 -15 -775
rect 24 -801 25 -761
rect 27 -801 28 -761
rect 253 -772 254 -747
rect 256 -772 257 -747
rect 261 -772 262 -747
rect 264 -772 265 -747
rect 291 -772 292 -747
rect 294 -772 295 -747
rect 335 -772 336 -747
rect 338 -772 339 -747
rect 380 -772 381 -747
rect 383 -772 384 -747
rect -52 -828 -51 -808
rect -49 -828 -48 -808
rect -68 -1106 -67 -1066
rect -65 -1106 -64 -1066
rect 2 -1101 3 -1081
rect 5 -1101 6 -1081
rect 45 -1107 46 -1067
rect 48 -1107 49 -1067
rect 274 -1078 275 -1053
rect 277 -1078 278 -1053
rect 282 -1078 283 -1053
rect 285 -1078 286 -1053
rect 312 -1078 313 -1053
rect 315 -1078 316 -1053
rect 356 -1078 357 -1053
rect 359 -1078 360 -1053
rect 401 -1078 402 -1053
rect 404 -1078 405 -1053
rect -31 -1134 -30 -1114
rect -28 -1134 -27 -1114
rect 339 -1318 340 -1293
rect 342 -1318 343 -1293
rect 347 -1318 348 -1293
rect 350 -1318 351 -1293
rect 377 -1318 378 -1293
rect 380 -1318 381 -1293
rect 421 -1318 422 -1293
rect 424 -1318 425 -1293
rect 466 -1318 467 -1293
rect 469 -1318 470 -1293
<< ndcontact >>
rect -390 -201 -386 -191
rect -382 -201 -378 -191
rect -354 -201 -350 -191
rect -346 -201 -342 -191
rect -338 -201 -334 -191
rect -310 -201 -306 -191
rect -302 -201 -298 -191
rect -294 -201 -290 -191
rect -259 -201 -255 -191
rect -251 -201 -247 -191
rect -70 -221 -66 -201
rect -62 -221 -58 -201
rect -107 -273 -103 -253
rect -99 -273 -95 -253
rect -37 -268 -33 -248
rect -29 -268 -25 -248
rect 231 -237 235 -227
rect 239 -237 243 -227
rect 267 -237 271 -227
rect 275 -237 279 -227
rect 283 -237 287 -227
rect 311 -237 315 -227
rect 319 -237 323 -227
rect 327 -237 331 -227
rect 362 -237 366 -227
rect 370 -237 374 -227
rect 6 -274 10 -254
rect 14 -274 18 -254
rect -80 -529 -76 -509
rect -72 -529 -68 -509
rect -117 -581 -113 -561
rect -109 -581 -105 -561
rect -47 -576 -43 -556
rect -39 -576 -35 -556
rect 221 -545 225 -535
rect 229 -545 233 -535
rect 257 -545 261 -535
rect 265 -545 269 -535
rect 273 -545 277 -535
rect 301 -545 305 -535
rect 309 -545 313 -535
rect 317 -545 321 -535
rect 352 -545 356 -535
rect 360 -545 364 -535
rect -4 -582 0 -562
rect 4 -582 8 -562
rect -56 -788 -52 -768
rect -48 -788 -44 -768
rect -93 -840 -89 -820
rect -85 -840 -81 -820
rect -23 -835 -19 -815
rect -15 -835 -11 -815
rect 245 -804 249 -794
rect 253 -804 257 -794
rect 281 -804 285 -794
rect 289 -804 293 -794
rect 297 -804 301 -794
rect 325 -804 329 -794
rect 333 -804 337 -794
rect 341 -804 345 -794
rect 376 -804 380 -794
rect 384 -804 388 -794
rect 20 -841 24 -821
rect 28 -841 32 -821
rect -35 -1094 -31 -1074
rect -27 -1094 -23 -1074
rect -72 -1146 -68 -1126
rect -64 -1146 -60 -1126
rect -2 -1141 2 -1121
rect 6 -1141 10 -1121
rect 266 -1110 270 -1100
rect 274 -1110 278 -1100
rect 302 -1110 306 -1100
rect 310 -1110 314 -1100
rect 318 -1110 322 -1100
rect 346 -1110 350 -1100
rect 354 -1110 358 -1100
rect 362 -1110 366 -1100
rect 397 -1110 401 -1100
rect 405 -1110 409 -1100
rect 41 -1147 45 -1127
rect 49 -1147 53 -1127
rect 331 -1350 335 -1340
rect 339 -1350 343 -1340
rect 367 -1350 371 -1340
rect 375 -1350 379 -1340
rect 383 -1350 387 -1340
rect 411 -1350 415 -1340
rect 419 -1350 423 -1340
rect 427 -1350 431 -1340
rect 462 -1350 466 -1340
rect 470 -1350 474 -1340
<< pdcontact >>
rect -386 -169 -382 -144
rect -378 -169 -374 -144
rect -370 -169 -366 -144
rect -348 -169 -344 -144
rect -340 -169 -336 -144
rect -304 -169 -300 -144
rect -296 -169 -292 -144
rect -259 -169 -255 -144
rect -251 -169 -247 -144
rect -107 -233 -103 -193
rect -99 -233 -95 -193
rect -37 -228 -33 -208
rect -29 -228 -25 -208
rect 6 -234 10 -194
rect 14 -234 18 -194
rect 235 -205 239 -180
rect 243 -205 247 -180
rect 251 -205 255 -180
rect 273 -205 277 -180
rect 281 -205 285 -180
rect 317 -205 321 -180
rect 325 -205 329 -180
rect 362 -205 366 -180
rect 370 -205 374 -180
rect -70 -261 -66 -241
rect -62 -261 -58 -241
rect -117 -541 -113 -501
rect -109 -541 -105 -501
rect -47 -536 -43 -516
rect -39 -536 -35 -516
rect -4 -542 0 -502
rect 4 -542 8 -502
rect 225 -513 229 -488
rect 233 -513 237 -488
rect 241 -513 245 -488
rect 263 -513 267 -488
rect 271 -513 275 -488
rect 307 -513 311 -488
rect 315 -513 319 -488
rect 352 -513 356 -488
rect 360 -513 364 -488
rect -80 -569 -76 -549
rect -72 -569 -68 -549
rect -93 -800 -89 -760
rect -85 -800 -81 -760
rect -23 -795 -19 -775
rect -15 -795 -11 -775
rect 20 -801 24 -761
rect 28 -801 32 -761
rect 249 -772 253 -747
rect 257 -772 261 -747
rect 265 -772 269 -747
rect 287 -772 291 -747
rect 295 -772 299 -747
rect 331 -772 335 -747
rect 339 -772 343 -747
rect 376 -772 380 -747
rect 384 -772 388 -747
rect -56 -828 -52 -808
rect -48 -828 -44 -808
rect -72 -1106 -68 -1066
rect -64 -1106 -60 -1066
rect -2 -1101 2 -1081
rect 6 -1101 10 -1081
rect 41 -1107 45 -1067
rect 49 -1107 53 -1067
rect 270 -1078 274 -1053
rect 278 -1078 282 -1053
rect 286 -1078 290 -1053
rect 308 -1078 312 -1053
rect 316 -1078 320 -1053
rect 352 -1078 356 -1053
rect 360 -1078 364 -1053
rect 397 -1078 401 -1053
rect 405 -1078 409 -1053
rect -35 -1134 -31 -1114
rect -27 -1134 -23 -1114
rect 335 -1318 339 -1293
rect 343 -1318 347 -1293
rect 351 -1318 355 -1293
rect 373 -1318 377 -1293
rect 381 -1318 385 -1293
rect 417 -1318 421 -1293
rect 425 -1318 429 -1293
rect 462 -1318 466 -1293
rect 470 -1318 474 -1293
<< polysilicon >>
rect -381 -144 -379 -141
rect -373 -144 -371 -141
rect -343 -144 -341 -141
rect -299 -144 -297 -141
rect -254 -144 -252 -141
rect -381 -176 -379 -169
rect -386 -180 -379 -176
rect -385 -191 -383 -180
rect -373 -188 -371 -169
rect -343 -177 -341 -169
rect -299 -177 -297 -169
rect -349 -179 -341 -177
rect -305 -179 -297 -177
rect -349 -191 -347 -179
rect -341 -191 -339 -182
rect -305 -191 -303 -179
rect -297 -191 -295 -182
rect -254 -191 -252 -169
rect 240 -180 242 -177
rect 248 -180 250 -177
rect 278 -180 280 -177
rect 322 -180 324 -177
rect 367 -180 369 -177
rect -102 -193 -100 -189
rect -385 -204 -383 -201
rect -349 -204 -347 -201
rect -341 -204 -339 -201
rect -305 -204 -303 -201
rect -297 -204 -295 -201
rect -254 -204 -252 -201
rect 11 -194 13 -190
rect -65 -201 -63 -194
rect -32 -208 -30 -194
rect -65 -224 -63 -221
rect -32 -231 -30 -228
rect -102 -253 -100 -233
rect 240 -212 242 -205
rect 235 -216 242 -212
rect 236 -227 238 -216
rect 248 -224 250 -205
rect 278 -213 280 -205
rect 322 -213 324 -205
rect 272 -215 280 -213
rect 316 -215 324 -213
rect 272 -227 274 -215
rect 280 -227 282 -218
rect 316 -227 318 -215
rect 324 -227 326 -218
rect 367 -227 369 -205
rect -65 -241 -63 -238
rect -32 -248 -30 -245
rect -102 -276 -100 -273
rect -65 -275 -63 -261
rect 11 -254 13 -234
rect 236 -240 238 -237
rect 272 -240 274 -237
rect 280 -240 282 -237
rect 316 -240 318 -237
rect 324 -240 326 -237
rect 367 -240 369 -237
rect -32 -275 -30 -268
rect 11 -277 13 -274
rect 230 -488 232 -485
rect 238 -488 240 -485
rect 268 -488 270 -485
rect 312 -488 314 -485
rect 357 -488 359 -485
rect -112 -501 -110 -497
rect 1 -502 3 -498
rect -75 -509 -73 -502
rect -42 -516 -40 -502
rect -75 -532 -73 -529
rect -42 -539 -40 -536
rect -112 -561 -110 -541
rect 230 -520 232 -513
rect 225 -524 232 -520
rect 226 -535 228 -524
rect 238 -532 240 -513
rect 268 -521 270 -513
rect 312 -521 314 -513
rect 262 -523 270 -521
rect 306 -523 314 -521
rect 262 -535 264 -523
rect 270 -535 272 -526
rect 306 -535 308 -523
rect 314 -535 316 -526
rect 357 -535 359 -513
rect -75 -549 -73 -546
rect -42 -556 -40 -553
rect -112 -584 -110 -581
rect -75 -583 -73 -569
rect 1 -562 3 -542
rect 226 -548 228 -545
rect 262 -548 264 -545
rect 270 -548 272 -545
rect 306 -548 308 -545
rect 314 -548 316 -545
rect 357 -548 359 -545
rect -42 -583 -40 -576
rect 1 -585 3 -582
rect 254 -747 256 -744
rect 262 -747 264 -744
rect 292 -747 294 -744
rect 336 -747 338 -744
rect 381 -747 383 -744
rect -88 -760 -86 -756
rect 25 -761 27 -757
rect -51 -768 -49 -761
rect -18 -775 -16 -761
rect -51 -791 -49 -788
rect -18 -798 -16 -795
rect -88 -820 -86 -800
rect 254 -779 256 -772
rect 249 -783 256 -779
rect 250 -794 252 -783
rect 262 -791 264 -772
rect 292 -780 294 -772
rect 336 -780 338 -772
rect 286 -782 294 -780
rect 330 -782 338 -780
rect 286 -794 288 -782
rect 294 -794 296 -785
rect 330 -794 332 -782
rect 338 -794 340 -785
rect 381 -794 383 -772
rect -51 -808 -49 -805
rect -18 -815 -16 -812
rect -88 -843 -86 -840
rect -51 -842 -49 -828
rect 25 -821 27 -801
rect 250 -807 252 -804
rect 286 -807 288 -804
rect 294 -807 296 -804
rect 330 -807 332 -804
rect 338 -807 340 -804
rect 381 -807 383 -804
rect -18 -842 -16 -835
rect 25 -844 27 -841
rect 275 -1053 277 -1050
rect 283 -1053 285 -1050
rect 313 -1053 315 -1050
rect 357 -1053 359 -1050
rect 402 -1053 404 -1050
rect -67 -1066 -65 -1062
rect 46 -1067 48 -1063
rect -30 -1074 -28 -1067
rect 3 -1081 5 -1067
rect -30 -1097 -28 -1094
rect 3 -1104 5 -1101
rect -67 -1126 -65 -1106
rect 275 -1085 277 -1078
rect 270 -1089 277 -1085
rect 271 -1100 273 -1089
rect 283 -1097 285 -1078
rect 313 -1086 315 -1078
rect 357 -1086 359 -1078
rect 307 -1088 315 -1086
rect 351 -1088 359 -1086
rect 307 -1100 309 -1088
rect 315 -1100 317 -1091
rect 351 -1100 353 -1088
rect 359 -1100 361 -1091
rect 402 -1100 404 -1078
rect -30 -1114 -28 -1111
rect 3 -1121 5 -1118
rect -67 -1149 -65 -1146
rect -30 -1148 -28 -1134
rect 46 -1127 48 -1107
rect 271 -1113 273 -1110
rect 307 -1113 309 -1110
rect 315 -1113 317 -1110
rect 351 -1113 353 -1110
rect 359 -1113 361 -1110
rect 402 -1113 404 -1110
rect 3 -1148 5 -1141
rect 46 -1150 48 -1147
rect 340 -1293 342 -1290
rect 348 -1293 350 -1290
rect 378 -1293 380 -1290
rect 422 -1293 424 -1290
rect 467 -1293 469 -1290
rect 340 -1325 342 -1318
rect 335 -1329 342 -1325
rect 336 -1340 338 -1329
rect 348 -1337 350 -1318
rect 378 -1326 380 -1318
rect 422 -1326 424 -1318
rect 372 -1328 380 -1326
rect 416 -1328 424 -1326
rect 372 -1340 374 -1328
rect 380 -1340 382 -1331
rect 416 -1340 418 -1328
rect 424 -1340 426 -1331
rect 467 -1340 469 -1318
rect 336 -1353 338 -1350
rect 372 -1353 374 -1350
rect 380 -1353 382 -1350
rect 416 -1353 418 -1350
rect 424 -1353 426 -1350
rect 467 -1353 469 -1350
<< polycontact >>
rect -390 -180 -386 -176
rect -377 -188 -373 -184
rect -354 -188 -349 -183
rect -339 -188 -334 -184
rect -310 -188 -305 -183
rect -258 -183 -254 -178
rect -295 -188 -290 -184
rect -66 -194 -62 -189
rect -33 -194 -29 -189
rect -106 -250 -102 -245
rect 231 -216 235 -212
rect 244 -224 248 -220
rect 267 -224 272 -219
rect 282 -224 287 -220
rect 311 -224 316 -219
rect 363 -219 367 -214
rect 326 -224 331 -220
rect 7 -251 11 -246
rect -66 -280 -62 -275
rect -33 -280 -29 -275
rect -76 -502 -72 -497
rect -43 -502 -39 -497
rect -116 -558 -112 -553
rect 221 -524 225 -520
rect 234 -532 238 -528
rect 257 -532 262 -527
rect 272 -532 277 -528
rect 301 -532 306 -527
rect 353 -527 357 -522
rect 316 -532 321 -528
rect -3 -559 1 -554
rect -76 -588 -72 -583
rect -43 -588 -39 -583
rect -52 -761 -48 -756
rect -19 -761 -15 -756
rect -92 -817 -88 -812
rect 245 -783 249 -779
rect 258 -791 262 -787
rect 281 -791 286 -786
rect 296 -791 301 -787
rect 325 -791 330 -786
rect 377 -786 381 -781
rect 340 -791 345 -787
rect 21 -818 25 -813
rect -52 -847 -48 -842
rect -19 -847 -15 -842
rect -31 -1067 -27 -1062
rect 2 -1067 6 -1062
rect -71 -1123 -67 -1118
rect 266 -1089 270 -1085
rect 279 -1097 283 -1093
rect 302 -1097 307 -1092
rect 317 -1097 322 -1093
rect 346 -1097 351 -1092
rect 398 -1092 402 -1087
rect 361 -1097 366 -1093
rect 42 -1124 46 -1119
rect -31 -1153 -27 -1148
rect 2 -1153 6 -1148
rect 331 -1329 335 -1325
rect 344 -1337 348 -1333
rect 367 -1337 372 -1332
rect 382 -1337 387 -1333
rect 411 -1337 416 -1332
rect 463 -1332 467 -1327
rect 426 -1337 431 -1333
<< metal1 >>
rect -392 -138 -239 -134
rect -386 -144 -382 -138
rect -348 -144 -344 -138
rect -304 -144 -300 -138
rect -259 -144 -255 -138
rect -336 -169 -323 -144
rect -292 -169 -279 -144
rect -135 -157 98 -152
rect -397 -180 -390 -176
rect -370 -177 -366 -169
rect -370 -180 -330 -177
rect -380 -188 -377 -184
rect -370 -191 -366 -180
rect -358 -188 -354 -183
rect -334 -188 -330 -180
rect -326 -183 -323 -169
rect -282 -178 -279 -169
rect -282 -183 -258 -178
rect -251 -179 -247 -169
rect -326 -188 -310 -183
rect -290 -188 -286 -184
rect -326 -191 -323 -188
rect -282 -191 -279 -183
rect -251 -184 -238 -179
rect -251 -191 -247 -184
rect -378 -201 -366 -191
rect -334 -201 -323 -191
rect -290 -201 -279 -191
rect -107 -193 -103 -157
rect -390 -206 -386 -201
rect -354 -206 -350 -201
rect -310 -206 -306 -201
rect -259 -206 -255 -201
rect -391 -210 -247 -206
rect -82 -225 -77 -170
rect -66 -189 -62 -182
rect -33 -189 -29 -182
rect 6 -194 10 -157
rect 53 -177 104 -171
rect 229 -174 382 -170
rect 26 -182 104 -177
rect 235 -180 239 -174
rect 273 -180 277 -174
rect 317 -180 321 -174
rect 362 -180 366 -174
rect -70 -225 -66 -221
rect -82 -229 -66 -225
rect -116 -250 -106 -245
rect -99 -246 -95 -233
rect -70 -241 -66 -229
rect -99 -251 -86 -246
rect -99 -253 -95 -251
rect -62 -226 -58 -221
rect -62 -230 -45 -226
rect -62 -241 -58 -230
rect -49 -240 -45 -230
rect -37 -240 -33 -228
rect -49 -245 -33 -240
rect -107 -312 -103 -273
rect -66 -293 -62 -280
rect -49 -303 -43 -245
rect -37 -248 -33 -245
rect -29 -241 -25 -228
rect 285 -205 298 -180
rect 329 -205 342 -180
rect 214 -216 231 -212
rect 251 -213 255 -205
rect 251 -216 291 -213
rect 241 -224 244 -220
rect 251 -227 255 -216
rect 263 -224 267 -219
rect 287 -224 291 -216
rect 295 -219 298 -205
rect 339 -214 342 -205
rect 339 -219 363 -214
rect 370 -215 374 -205
rect 295 -224 311 -219
rect 331 -224 335 -220
rect 295 -227 298 -224
rect 339 -227 342 -219
rect 370 -220 383 -215
rect 370 -227 374 -220
rect -29 -245 -8 -241
rect -29 -248 -25 -245
rect -14 -246 -8 -245
rect -14 -251 -4 -246
rect 2 -251 7 -246
rect 14 -247 18 -234
rect 243 -237 255 -227
rect 287 -237 298 -227
rect 331 -237 342 -227
rect 231 -242 235 -237
rect 267 -242 271 -237
rect 311 -242 315 -237
rect 362 -242 366 -237
rect 230 -246 374 -242
rect 14 -252 31 -247
rect 14 -254 18 -252
rect 56 -255 74 -249
rect -33 -293 -29 -280
rect 6 -312 10 -274
rect 56 -292 64 -255
rect -135 -320 74 -312
rect -145 -465 88 -460
rect -117 -501 -113 -465
rect -92 -533 -87 -478
rect -76 -497 -72 -490
rect -43 -497 -39 -490
rect -4 -502 0 -465
rect 43 -485 94 -479
rect 219 -482 372 -478
rect 16 -490 94 -485
rect 225 -488 229 -482
rect 263 -488 267 -482
rect 307 -488 311 -482
rect 352 -488 356 -482
rect -80 -533 -76 -529
rect -92 -537 -76 -533
rect -126 -558 -116 -553
rect -109 -554 -105 -541
rect -80 -549 -76 -537
rect -109 -559 -96 -554
rect -109 -561 -105 -559
rect -72 -534 -68 -529
rect -72 -538 -55 -534
rect -72 -549 -68 -538
rect -59 -548 -55 -538
rect -47 -548 -43 -536
rect -59 -553 -43 -548
rect -117 -620 -113 -581
rect -76 -601 -72 -588
rect -59 -611 -53 -553
rect -47 -556 -43 -553
rect -39 -549 -35 -536
rect 275 -513 288 -488
rect 319 -513 332 -488
rect 204 -524 221 -520
rect 241 -521 245 -513
rect 241 -524 281 -521
rect 231 -532 234 -528
rect 241 -535 245 -524
rect 253 -532 257 -527
rect 277 -532 281 -524
rect 285 -527 288 -513
rect 329 -522 332 -513
rect 329 -527 353 -522
rect 360 -523 364 -513
rect 285 -532 301 -527
rect 321 -532 325 -528
rect 285 -535 288 -532
rect 329 -535 332 -527
rect 360 -528 373 -523
rect 360 -535 364 -528
rect -39 -553 -18 -549
rect -39 -556 -35 -553
rect -24 -554 -18 -553
rect -24 -559 -14 -554
rect -8 -559 -3 -554
rect 4 -555 8 -542
rect 233 -545 245 -535
rect 277 -545 288 -535
rect 321 -545 332 -535
rect 221 -550 225 -545
rect 257 -550 261 -545
rect 301 -550 305 -545
rect 352 -550 356 -545
rect 220 -554 364 -550
rect 4 -560 21 -555
rect 4 -562 8 -560
rect 46 -563 64 -557
rect -43 -601 -39 -588
rect -4 -620 0 -582
rect 46 -600 54 -563
rect -145 -628 64 -620
rect -121 -724 112 -719
rect -93 -760 -89 -724
rect -68 -792 -63 -737
rect -52 -756 -48 -749
rect -19 -756 -15 -749
rect 20 -761 24 -724
rect 67 -744 118 -738
rect 243 -741 396 -737
rect 40 -749 118 -744
rect 249 -747 253 -741
rect 287 -747 291 -741
rect 331 -747 335 -741
rect 376 -747 380 -741
rect -56 -792 -52 -788
rect -68 -796 -52 -792
rect -102 -817 -92 -812
rect -85 -813 -81 -800
rect -56 -808 -52 -796
rect -85 -818 -72 -813
rect -85 -820 -81 -818
rect -48 -793 -44 -788
rect -48 -797 -31 -793
rect -48 -808 -44 -797
rect -35 -807 -31 -797
rect -23 -807 -19 -795
rect -35 -812 -19 -807
rect -93 -879 -89 -840
rect -52 -860 -48 -847
rect -35 -870 -29 -812
rect -23 -815 -19 -812
rect -15 -808 -11 -795
rect 299 -772 312 -747
rect 343 -772 356 -747
rect 228 -783 245 -779
rect 265 -780 269 -772
rect 265 -783 305 -780
rect 255 -791 258 -787
rect 265 -794 269 -783
rect 277 -791 281 -786
rect 301 -791 305 -783
rect 309 -786 312 -772
rect 353 -781 356 -772
rect 353 -786 377 -781
rect 384 -782 388 -772
rect 309 -791 325 -786
rect 345 -791 349 -787
rect 309 -794 312 -791
rect 353 -794 356 -786
rect 384 -787 397 -782
rect 384 -794 388 -787
rect -15 -812 6 -808
rect -15 -815 -11 -812
rect 0 -813 6 -812
rect 0 -818 10 -813
rect 16 -818 21 -813
rect 28 -814 32 -801
rect 257 -804 269 -794
rect 301 -804 312 -794
rect 345 -804 356 -794
rect 245 -809 249 -804
rect 281 -809 285 -804
rect 325 -809 329 -804
rect 376 -809 380 -804
rect 244 -813 388 -809
rect 28 -819 45 -814
rect 28 -821 32 -819
rect 70 -822 88 -816
rect -19 -860 -15 -847
rect 20 -879 24 -841
rect 70 -859 78 -822
rect -121 -887 88 -879
rect -100 -1030 133 -1025
rect -72 -1066 -68 -1030
rect -47 -1098 -42 -1043
rect -31 -1062 -27 -1055
rect 2 -1062 6 -1055
rect 41 -1067 45 -1030
rect 88 -1050 139 -1044
rect 264 -1047 417 -1043
rect 61 -1055 139 -1050
rect 270 -1053 274 -1047
rect 308 -1053 312 -1047
rect 352 -1053 356 -1047
rect 397 -1053 401 -1047
rect -35 -1098 -31 -1094
rect -47 -1102 -31 -1098
rect -81 -1123 -71 -1118
rect -64 -1119 -60 -1106
rect -35 -1114 -31 -1102
rect -64 -1124 -51 -1119
rect -64 -1126 -60 -1124
rect -27 -1099 -23 -1094
rect -27 -1103 -10 -1099
rect -27 -1114 -23 -1103
rect -14 -1113 -10 -1103
rect -2 -1113 2 -1101
rect -14 -1118 2 -1113
rect -72 -1185 -68 -1146
rect -31 -1166 -27 -1153
rect -14 -1176 -8 -1118
rect -2 -1121 2 -1118
rect 6 -1114 10 -1101
rect 320 -1078 333 -1053
rect 364 -1078 377 -1053
rect 249 -1089 266 -1085
rect 286 -1086 290 -1078
rect 286 -1089 326 -1086
rect 276 -1097 279 -1093
rect 286 -1100 290 -1089
rect 298 -1097 302 -1092
rect 322 -1097 326 -1089
rect 330 -1092 333 -1078
rect 374 -1087 377 -1078
rect 374 -1092 398 -1087
rect 405 -1088 409 -1078
rect 330 -1097 346 -1092
rect 366 -1097 370 -1093
rect 330 -1100 333 -1097
rect 374 -1100 377 -1092
rect 405 -1093 418 -1088
rect 405 -1100 409 -1093
rect 6 -1118 27 -1114
rect 6 -1121 10 -1118
rect 21 -1119 27 -1118
rect 21 -1124 31 -1119
rect 37 -1124 42 -1119
rect 49 -1120 53 -1107
rect 278 -1110 290 -1100
rect 322 -1110 333 -1100
rect 366 -1110 377 -1100
rect 266 -1115 270 -1110
rect 302 -1115 306 -1110
rect 346 -1115 350 -1110
rect 397 -1115 401 -1110
rect 265 -1119 409 -1115
rect 49 -1125 66 -1120
rect 49 -1127 53 -1125
rect 91 -1128 109 -1122
rect 2 -1166 6 -1153
rect 41 -1185 45 -1147
rect 91 -1165 99 -1128
rect -100 -1193 109 -1185
rect 329 -1287 482 -1283
rect 335 -1293 339 -1287
rect 373 -1293 377 -1287
rect 417 -1293 421 -1287
rect 462 -1293 466 -1287
rect 385 -1318 398 -1293
rect 429 -1318 442 -1293
rect 324 -1329 331 -1325
rect 351 -1326 355 -1318
rect 351 -1329 391 -1326
rect 341 -1337 344 -1333
rect 351 -1340 355 -1329
rect 363 -1337 367 -1332
rect 387 -1337 391 -1329
rect 395 -1332 398 -1318
rect 439 -1327 442 -1318
rect 439 -1332 463 -1327
rect 470 -1328 474 -1318
rect 395 -1337 411 -1332
rect 431 -1337 435 -1333
rect 395 -1340 398 -1337
rect 439 -1340 442 -1332
rect 470 -1333 483 -1328
rect 470 -1340 474 -1333
rect 343 -1350 355 -1340
rect 387 -1350 398 -1340
rect 431 -1350 442 -1340
rect 331 -1355 335 -1350
rect 367 -1355 371 -1350
rect 411 -1355 415 -1350
rect 462 -1355 466 -1350
rect 330 -1359 474 -1355
<< m2contact >>
rect -82 -170 -76 -165
rect -66 -182 -61 -177
rect -34 -182 -29 -177
rect 18 -182 26 -177
rect -121 -250 -116 -245
rect -86 -251 -80 -246
rect -66 -298 -61 -293
rect 209 -217 214 -212
rect -4 -251 2 -246
rect 31 -252 37 -247
rect -33 -298 -28 -293
rect -49 -309 -43 -303
rect 56 -298 64 -292
rect -92 -478 -86 -473
rect -76 -490 -71 -485
rect -44 -490 -39 -485
rect 8 -490 16 -485
rect -131 -558 -126 -553
rect -96 -559 -90 -554
rect -76 -606 -71 -601
rect 199 -525 204 -520
rect -14 -559 -8 -554
rect 21 -560 27 -555
rect -43 -606 -38 -601
rect -59 -617 -53 -611
rect 46 -606 54 -600
rect -68 -737 -62 -732
rect -52 -749 -47 -744
rect -20 -749 -15 -744
rect 32 -749 40 -744
rect -107 -817 -102 -812
rect -72 -818 -66 -813
rect -52 -865 -47 -860
rect 223 -784 228 -779
rect 10 -818 16 -813
rect 45 -819 51 -814
rect -19 -865 -14 -860
rect -35 -876 -29 -870
rect 70 -865 78 -859
rect -47 -1043 -41 -1038
rect -31 -1055 -26 -1050
rect 1 -1055 6 -1050
rect 53 -1055 61 -1050
rect -86 -1123 -81 -1118
rect -51 -1124 -45 -1119
rect -31 -1171 -26 -1166
rect 244 -1090 249 -1085
rect 31 -1124 37 -1119
rect 66 -1125 72 -1120
rect 2 -1171 7 -1166
rect -14 -1182 -8 -1176
rect 91 -1171 99 -1165
<< metal2 >>
rect -76 -170 37 -165
rect -121 -182 -66 -177
rect -61 -182 -34 -177
rect -29 -182 18 -177
rect -121 -245 -117 -182
rect -86 -293 -80 -251
rect -4 -292 2 -251
rect 31 -247 37 -170
rect -87 -298 -66 -293
rect -61 -298 -33 -293
rect -28 -298 -14 -293
rect -4 -298 56 -292
rect 209 -305 214 -217
rect -43 -309 214 -305
rect -86 -478 27 -473
rect -131 -490 -76 -485
rect -71 -490 -44 -485
rect -39 -490 8 -485
rect -131 -553 -127 -490
rect -96 -601 -90 -559
rect -14 -600 -8 -559
rect 21 -555 27 -478
rect -97 -606 -76 -601
rect -71 -606 -43 -601
rect -38 -606 -24 -601
rect -14 -606 46 -600
rect 199 -613 204 -525
rect -53 -617 204 -613
rect -62 -737 51 -732
rect -107 -749 -52 -744
rect -47 -749 -20 -744
rect -15 -749 32 -744
rect -107 -812 -103 -749
rect -72 -860 -66 -818
rect 10 -859 16 -818
rect 45 -814 51 -737
rect -73 -865 -52 -860
rect -47 -865 -19 -860
rect -14 -865 0 -860
rect 10 -865 70 -859
rect 223 -872 228 -784
rect -29 -876 228 -872
rect -41 -1043 72 -1038
rect -86 -1055 -31 -1050
rect -26 -1055 1 -1050
rect 6 -1055 53 -1050
rect -86 -1118 -82 -1055
rect -51 -1166 -45 -1124
rect 31 -1165 37 -1124
rect 66 -1120 72 -1043
rect -52 -1171 -31 -1166
rect -26 -1171 2 -1166
rect 7 -1171 21 -1166
rect 31 -1171 91 -1165
rect 244 -1178 249 -1090
rect -8 -1182 249 -1178
<< labels >>
rlabel metal1 -50 -319 64 -313 1 GND
rlabel metal1 -26 -157 88 -152 5 VDD
rlabel metal1 56 -255 72 -249 1 p0
rlabel metal1 332 -223 334 -221 1 clk
rlabel metal1 264 -223 265 -221 1 clk
rlabel metal1 245 -172 247 -171 5 vdd
rlabel metal1 239 -244 242 -243 1 gnd
rlabel metal1 241 -223 243 -221 1 clk
rlabel metal1 376 -218 379 -216 1 s0_reg
rlabel metal1 226 -215 228 -213 1 s0
rlabel metal1 -49 -302 -43 -298 1 s0
rlabel metal1 -60 -627 54 -621 1 GND
rlabel metal1 -36 -465 78 -460 5 VDD
rlabel metal1 322 -531 324 -529 1 clk
rlabel metal1 254 -531 255 -529 1 clk
rlabel metal1 235 -480 237 -479 5 vdd
rlabel metal1 229 -552 232 -551 1 gnd
rlabel metal1 231 -531 233 -529 1 clk
rlabel metal1 -36 -886 78 -880 1 GND
rlabel metal1 -12 -724 102 -719 5 VDD
rlabel metal1 346 -790 348 -788 1 clk
rlabel metal1 278 -790 279 -788 1 clk
rlabel metal1 259 -739 261 -738 5 vdd
rlabel metal1 253 -811 256 -810 1 gnd
rlabel metal1 255 -790 257 -788 1 clk
rlabel metal1 341 -1336 343 -1334 1 clk
rlabel metal1 339 -1357 342 -1356 1 gnd
rlabel metal1 345 -1285 347 -1284 5 vdd
rlabel metal1 364 -1336 365 -1334 1 clk
rlabel metal1 432 -1336 434 -1334 1 clk
rlabel metal1 326 -1328 328 -1326 1 out_carry
rlabel metal1 475 -1331 480 -1329 1 out_carry_reg
rlabel metal1 -15 -1192 99 -1186 1 GND
rlabel metal1 9 -1030 123 -1025 5 VDD
rlabel metal1 367 -1096 369 -1094 1 clk
rlabel metal1 299 -1096 300 -1094 1 clk
rlabel metal1 280 -1045 282 -1044 5 vdd
rlabel metal1 274 -1117 277 -1116 1 gnd
rlabel metal1 276 -1096 278 -1094 1 clk
rlabel metal1 216 -523 218 -521 1 s1
rlabel metal1 366 -526 369 -524 1 s1_reg
rlabel metal1 -59 -610 -53 -606 1 s1
rlabel metal1 -35 -869 -29 -865 1 s2
rlabel metal1 -14 -1175 -8 -1171 1 s3
rlabel metal1 240 -782 242 -780 1 s2
rlabel metal1 390 -785 393 -783 1 s2_reg
rlabel metal1 411 -1091 414 -1089 1 s3_reg
rlabel metal1 261 -1088 263 -1086 1 s3
rlabel metal1 52 -484 89 -479 1 c0
rlabel metal1 46 -563 62 -557 1 p1
rlabel metal1 70 -822 86 -816 1 p2
rlabel metal1 76 -743 113 -738 1 c1
rlabel metal1 91 -1128 107 -1122 1 p3
rlabel metal1 97 -1049 134 -1044 1 c2
rlabel metal1 62 -176 99 -171 1 carry_reg
rlabel metal1 -380 -187 -378 -185 1 clk
rlabel metal1 -382 -208 -379 -207 1 gnd
rlabel metal1 -376 -136 -374 -135 5 vdd
rlabel metal1 -357 -187 -356 -185 1 clk
rlabel metal1 -289 -187 -287 -185 1 clk
rlabel metal1 -246 -182 -241 -180 1 carry_reg
rlabel metal1 -395 -179 -393 -177 3 carry
<< end >>
