magic
tech scmos
timestamp 1732067555
<< nwell >>
rect -82 -2340 -50 -2303
rect -44 -2340 -18 -2303
rect 0 -2340 26 -2303
rect 45 -2340 71 -2303
rect 184 -2447 218 -2411
rect 225 -2448 249 -2424
rect 482 -2430 507 -2373
rect 519 -2458 544 -2418
rect 552 -2425 577 -2385
rect 595 -2431 620 -2374
rect 824 -2398 856 -2361
rect 862 -2398 888 -2361
rect 906 -2398 932 -2361
rect 951 -2398 977 -2361
rect 85 -2488 119 -2464
rect 125 -2489 149 -2465
rect -845 -2549 -813 -2512
rect -807 -2549 -781 -2512
rect -763 -2549 -737 -2512
rect -718 -2549 -692 -2512
rect -632 -2549 -600 -2512
rect -594 -2549 -568 -2512
rect -550 -2549 -524 -2512
rect -505 -2549 -479 -2512
rect -385 -2599 -360 -2542
rect -348 -2627 -323 -2587
rect -315 -2594 -290 -2554
rect -272 -2600 -247 -2543
rect -139 -2556 -105 -2532
rect -99 -2557 -75 -2533
rect 92 -2731 126 -2707
rect 132 -2732 156 -2708
rect 472 -2738 497 -2681
rect 194 -2812 228 -2776
rect 345 -2783 379 -2747
rect 386 -2784 410 -2760
rect 509 -2766 534 -2726
rect 542 -2733 567 -2693
rect 585 -2739 610 -2682
rect 814 -2706 846 -2669
rect 852 -2706 878 -2669
rect 896 -2706 922 -2669
rect 941 -2706 967 -2669
rect 235 -2813 259 -2789
rect -830 -2878 -798 -2841
rect -792 -2878 -766 -2841
rect -748 -2878 -722 -2841
rect -703 -2878 -677 -2841
rect -617 -2878 -585 -2841
rect -579 -2878 -553 -2841
rect -535 -2878 -509 -2841
rect -490 -2878 -464 -2841
rect 95 -2853 129 -2829
rect 135 -2854 159 -2830
rect -370 -2928 -345 -2871
rect -333 -2956 -308 -2916
rect -300 -2923 -275 -2883
rect -257 -2929 -232 -2872
rect -124 -2885 -90 -2861
rect -84 -2886 -60 -2862
rect 90 -2995 124 -2971
rect 130 -2996 154 -2972
rect 496 -2997 521 -2940
rect 533 -3025 558 -2985
rect 566 -2992 591 -2952
rect 609 -2998 634 -2941
rect 838 -2965 870 -2928
rect 876 -2965 902 -2928
rect 920 -2965 946 -2928
rect 965 -2965 991 -2928
rect 192 -3076 226 -3040
rect 233 -3077 257 -3053
rect -806 -3145 -774 -3108
rect -768 -3145 -742 -3108
rect -724 -3145 -698 -3108
rect -679 -3145 -653 -3108
rect -593 -3145 -561 -3108
rect -555 -3145 -529 -3108
rect -511 -3145 -485 -3108
rect -466 -3145 -440 -3108
rect 93 -3117 127 -3093
rect 133 -3118 157 -3094
rect 301 -3103 335 -3067
rect 342 -3104 366 -3080
rect -346 -3195 -321 -3138
rect -309 -3223 -284 -3183
rect -276 -3190 -251 -3150
rect -233 -3196 -208 -3139
rect -100 -3152 -66 -3128
rect -60 -3153 -36 -3129
rect 194 -3163 228 -3127
rect 235 -3164 259 -3140
rect 100 -3196 134 -3172
rect 140 -3197 164 -3173
rect 517 -3303 542 -3246
rect 96 -3340 130 -3316
rect 136 -3341 160 -3317
rect 554 -3331 579 -3291
rect 587 -3298 612 -3258
rect 630 -3304 655 -3247
rect 859 -3271 891 -3234
rect 897 -3271 923 -3234
rect 941 -3271 967 -3234
rect 986 -3271 1012 -3234
rect -777 -3455 -745 -3418
rect -739 -3455 -713 -3418
rect -695 -3455 -669 -3418
rect -650 -3455 -624 -3418
rect -564 -3455 -532 -3418
rect -526 -3455 -500 -3418
rect -482 -3455 -456 -3418
rect -437 -3455 -411 -3418
rect 198 -3421 232 -3385
rect 239 -3422 263 -3398
rect -317 -3505 -292 -3448
rect -280 -3533 -255 -3493
rect -247 -3500 -222 -3460
rect -204 -3506 -179 -3449
rect -71 -3462 -37 -3438
rect -31 -3463 -7 -3439
rect 99 -3462 133 -3438
rect 139 -3463 163 -3439
rect 307 -3448 341 -3412
rect 348 -3449 372 -3425
rect 409 -3472 443 -3436
rect 200 -3508 234 -3472
rect 450 -3473 474 -3449
rect 599 -3473 631 -3436
rect 637 -3473 663 -3436
rect 681 -3473 707 -3436
rect 726 -3473 752 -3436
rect 241 -3509 265 -3485
rect 106 -3541 140 -3517
rect 146 -3542 170 -3518
rect 106 -3623 140 -3599
rect 146 -3624 170 -3600
<< ntransistor >>
rect -75 -2366 -73 -2356
rect -39 -2366 -37 -2356
rect -31 -2366 -29 -2356
rect 5 -2366 7 -2356
rect 13 -2366 15 -2356
rect 56 -2366 58 -2356
rect 530 -2408 532 -2388
rect 236 -2462 238 -2456
rect 493 -2460 495 -2440
rect 195 -2468 197 -2462
rect 205 -2468 207 -2462
rect 563 -2455 565 -2435
rect 831 -2424 833 -2414
rect 867 -2424 869 -2414
rect 875 -2424 877 -2414
rect 911 -2424 913 -2414
rect 919 -2424 921 -2414
rect 962 -2424 964 -2414
rect 606 -2461 608 -2441
rect 96 -2514 98 -2502
rect 106 -2514 108 -2502
rect 136 -2503 138 -2497
rect -838 -2575 -836 -2565
rect -802 -2575 -800 -2565
rect -794 -2575 -792 -2565
rect -758 -2575 -756 -2565
rect -750 -2575 -748 -2565
rect -707 -2575 -705 -2565
rect -625 -2575 -623 -2565
rect -589 -2575 -587 -2565
rect -581 -2575 -579 -2565
rect -545 -2575 -543 -2565
rect -537 -2575 -535 -2565
rect -494 -2575 -492 -2565
rect -337 -2577 -335 -2557
rect -128 -2582 -126 -2570
rect -118 -2582 -116 -2570
rect -88 -2571 -86 -2565
rect -374 -2629 -372 -2609
rect -304 -2624 -302 -2604
rect -261 -2630 -259 -2610
rect 520 -2716 522 -2696
rect 103 -2757 105 -2745
rect 113 -2757 115 -2745
rect 143 -2746 145 -2740
rect 483 -2768 485 -2748
rect 553 -2763 555 -2743
rect 821 -2732 823 -2722
rect 857 -2732 859 -2722
rect 865 -2732 867 -2722
rect 901 -2732 903 -2722
rect 909 -2732 911 -2722
rect 952 -2732 954 -2722
rect 596 -2769 598 -2749
rect 397 -2798 399 -2792
rect 356 -2804 358 -2798
rect 366 -2804 368 -2798
rect 246 -2827 248 -2821
rect 205 -2833 207 -2827
rect 215 -2833 217 -2827
rect -823 -2904 -821 -2894
rect -787 -2904 -785 -2894
rect -779 -2904 -777 -2894
rect -743 -2904 -741 -2894
rect -735 -2904 -733 -2894
rect -692 -2904 -690 -2894
rect -610 -2904 -608 -2894
rect -574 -2904 -572 -2894
rect -566 -2904 -564 -2894
rect -530 -2904 -528 -2894
rect -522 -2904 -520 -2894
rect -479 -2904 -477 -2894
rect -322 -2906 -320 -2886
rect 106 -2879 108 -2867
rect 116 -2879 118 -2867
rect 146 -2868 148 -2862
rect -113 -2911 -111 -2899
rect -103 -2911 -101 -2899
rect -73 -2900 -71 -2894
rect -359 -2958 -357 -2938
rect -289 -2953 -287 -2933
rect -246 -2959 -244 -2939
rect 544 -2975 546 -2955
rect 101 -3021 103 -3009
rect 111 -3021 113 -3009
rect 141 -3010 143 -3004
rect 507 -3027 509 -3007
rect 577 -3022 579 -3002
rect 845 -2991 847 -2981
rect 881 -2991 883 -2981
rect 889 -2991 891 -2981
rect 925 -2991 927 -2981
rect 933 -2991 935 -2981
rect 976 -2991 978 -2981
rect 620 -3028 622 -3008
rect 244 -3091 246 -3085
rect 203 -3097 205 -3091
rect 213 -3097 215 -3091
rect 353 -3118 355 -3112
rect 312 -3124 314 -3118
rect 322 -3124 324 -3118
rect -799 -3171 -797 -3161
rect -763 -3171 -761 -3161
rect -755 -3171 -753 -3161
rect -719 -3171 -717 -3161
rect -711 -3171 -709 -3161
rect -668 -3171 -666 -3161
rect -586 -3171 -584 -3161
rect -550 -3171 -548 -3161
rect -542 -3171 -540 -3161
rect -506 -3171 -504 -3161
rect -498 -3171 -496 -3161
rect -455 -3171 -453 -3161
rect -298 -3173 -296 -3153
rect 104 -3143 106 -3131
rect 114 -3143 116 -3131
rect 144 -3132 146 -3126
rect -89 -3178 -87 -3166
rect -79 -3178 -77 -3166
rect -49 -3167 -47 -3161
rect -335 -3225 -333 -3205
rect -265 -3220 -263 -3200
rect 246 -3178 248 -3172
rect -222 -3226 -220 -3206
rect 205 -3184 207 -3178
rect 215 -3184 217 -3178
rect 111 -3222 113 -3210
rect 121 -3222 123 -3210
rect 151 -3211 153 -3205
rect 565 -3281 567 -3261
rect 528 -3333 530 -3313
rect 598 -3328 600 -3308
rect 866 -3297 868 -3287
rect 902 -3297 904 -3287
rect 910 -3297 912 -3287
rect 946 -3297 948 -3287
rect 954 -3297 956 -3287
rect 997 -3297 999 -3287
rect 641 -3334 643 -3314
rect 107 -3366 109 -3354
rect 117 -3366 119 -3354
rect 147 -3355 149 -3349
rect 250 -3436 252 -3430
rect -770 -3481 -768 -3471
rect -734 -3481 -732 -3471
rect -726 -3481 -724 -3471
rect -690 -3481 -688 -3471
rect -682 -3481 -680 -3471
rect -639 -3481 -637 -3471
rect -557 -3481 -555 -3471
rect -521 -3481 -519 -3471
rect -513 -3481 -511 -3471
rect -477 -3481 -475 -3471
rect -469 -3481 -467 -3471
rect -426 -3481 -424 -3471
rect 209 -3442 211 -3436
rect 219 -3442 221 -3436
rect -269 -3483 -267 -3463
rect -60 -3488 -58 -3476
rect -50 -3488 -48 -3476
rect -20 -3477 -18 -3471
rect 359 -3463 361 -3457
rect 318 -3469 320 -3463
rect 328 -3469 330 -3463
rect 110 -3488 112 -3476
rect 120 -3488 122 -3476
rect 150 -3477 152 -3471
rect -306 -3535 -304 -3515
rect -236 -3530 -234 -3510
rect 461 -3487 463 -3481
rect -193 -3536 -191 -3516
rect 420 -3493 422 -3487
rect 430 -3493 432 -3487
rect 606 -3499 608 -3489
rect 642 -3499 644 -3489
rect 650 -3499 652 -3489
rect 686 -3499 688 -3489
rect 694 -3499 696 -3489
rect 737 -3499 739 -3489
rect 252 -3523 254 -3517
rect 211 -3529 213 -3523
rect 221 -3529 223 -3523
rect 117 -3567 119 -3555
rect 127 -3567 129 -3555
rect 157 -3556 159 -3550
rect 117 -3649 119 -3637
rect 127 -3649 129 -3637
rect 157 -3638 159 -3632
<< ptransistor >>
rect -71 -2334 -69 -2309
rect -63 -2334 -61 -2309
rect -33 -2334 -31 -2309
rect 11 -2334 13 -2309
rect 56 -2334 58 -2309
rect 195 -2441 197 -2417
rect 205 -2441 207 -2417
rect 493 -2420 495 -2380
rect 563 -2415 565 -2395
rect 236 -2442 238 -2430
rect 606 -2421 608 -2381
rect 835 -2392 837 -2367
rect 843 -2392 845 -2367
rect 873 -2392 875 -2367
rect 917 -2392 919 -2367
rect 962 -2392 964 -2367
rect 530 -2448 532 -2428
rect 96 -2482 98 -2470
rect 106 -2482 108 -2470
rect 136 -2483 138 -2471
rect -834 -2543 -832 -2518
rect -826 -2543 -824 -2518
rect -796 -2543 -794 -2518
rect -752 -2543 -750 -2518
rect -707 -2543 -705 -2518
rect -621 -2543 -619 -2518
rect -613 -2543 -611 -2518
rect -583 -2543 -581 -2518
rect -539 -2543 -537 -2518
rect -494 -2543 -492 -2518
rect -374 -2589 -372 -2549
rect -128 -2550 -126 -2538
rect -118 -2550 -116 -2538
rect -304 -2584 -302 -2564
rect -261 -2590 -259 -2550
rect -88 -2551 -86 -2539
rect -337 -2617 -335 -2597
rect 103 -2725 105 -2713
rect 113 -2725 115 -2713
rect 143 -2726 145 -2714
rect 483 -2728 485 -2688
rect 553 -2723 555 -2703
rect 596 -2729 598 -2689
rect 825 -2700 827 -2675
rect 833 -2700 835 -2675
rect 863 -2700 865 -2675
rect 907 -2700 909 -2675
rect 952 -2700 954 -2675
rect 356 -2777 358 -2753
rect 366 -2777 368 -2753
rect 205 -2806 207 -2782
rect 215 -2806 217 -2782
rect 246 -2807 248 -2795
rect 397 -2778 399 -2766
rect 520 -2756 522 -2736
rect 106 -2847 108 -2835
rect 116 -2847 118 -2835
rect -819 -2872 -817 -2847
rect -811 -2872 -809 -2847
rect -781 -2872 -779 -2847
rect -737 -2872 -735 -2847
rect -692 -2872 -690 -2847
rect -606 -2872 -604 -2847
rect -598 -2872 -596 -2847
rect -568 -2872 -566 -2847
rect -524 -2872 -522 -2847
rect -479 -2872 -477 -2847
rect -359 -2918 -357 -2878
rect -113 -2879 -111 -2867
rect -103 -2879 -101 -2867
rect 146 -2848 148 -2836
rect -289 -2913 -287 -2893
rect -246 -2919 -244 -2879
rect -73 -2880 -71 -2868
rect -322 -2946 -320 -2926
rect 101 -2989 103 -2977
rect 111 -2989 113 -2977
rect 141 -2990 143 -2978
rect 507 -2987 509 -2947
rect 577 -2982 579 -2962
rect 620 -2988 622 -2948
rect 849 -2959 851 -2934
rect 857 -2959 859 -2934
rect 887 -2959 889 -2934
rect 931 -2959 933 -2934
rect 976 -2959 978 -2934
rect 544 -3015 546 -2995
rect 203 -3070 205 -3046
rect 213 -3070 215 -3046
rect 244 -3071 246 -3059
rect 312 -3097 314 -3073
rect 322 -3097 324 -3073
rect 104 -3111 106 -3099
rect 114 -3111 116 -3099
rect -795 -3139 -793 -3114
rect -787 -3139 -785 -3114
rect -757 -3139 -755 -3114
rect -713 -3139 -711 -3114
rect -668 -3139 -666 -3114
rect -582 -3139 -580 -3114
rect -574 -3139 -572 -3114
rect -544 -3139 -542 -3114
rect -500 -3139 -498 -3114
rect -455 -3139 -453 -3114
rect 144 -3112 146 -3100
rect 353 -3098 355 -3086
rect -335 -3185 -333 -3145
rect -89 -3146 -87 -3134
rect -79 -3146 -77 -3134
rect -265 -3180 -263 -3160
rect -222 -3186 -220 -3146
rect -49 -3147 -47 -3135
rect 205 -3157 207 -3133
rect 215 -3157 217 -3133
rect -298 -3213 -296 -3193
rect 111 -3190 113 -3178
rect 121 -3190 123 -3178
rect 246 -3158 248 -3146
rect 151 -3191 153 -3179
rect 528 -3293 530 -3253
rect 598 -3288 600 -3268
rect 641 -3294 643 -3254
rect 870 -3265 872 -3240
rect 878 -3265 880 -3240
rect 908 -3265 910 -3240
rect 952 -3265 954 -3240
rect 997 -3265 999 -3240
rect 107 -3334 109 -3322
rect 117 -3334 119 -3322
rect 147 -3335 149 -3323
rect 565 -3321 567 -3301
rect 209 -3415 211 -3391
rect 219 -3415 221 -3391
rect -766 -3449 -764 -3424
rect -758 -3449 -756 -3424
rect -728 -3449 -726 -3424
rect -684 -3449 -682 -3424
rect -639 -3449 -637 -3424
rect -553 -3449 -551 -3424
rect -545 -3449 -543 -3424
rect -515 -3449 -513 -3424
rect -471 -3449 -469 -3424
rect -426 -3449 -424 -3424
rect 250 -3416 252 -3404
rect -306 -3495 -304 -3455
rect -60 -3456 -58 -3444
rect -50 -3456 -48 -3444
rect 318 -3442 320 -3418
rect 328 -3442 330 -3418
rect -236 -3490 -234 -3470
rect -193 -3496 -191 -3456
rect -20 -3457 -18 -3445
rect 110 -3456 112 -3444
rect 120 -3456 122 -3444
rect 150 -3457 152 -3445
rect 359 -3443 361 -3431
rect 420 -3466 422 -3442
rect 430 -3466 432 -3442
rect -269 -3523 -267 -3503
rect 211 -3502 213 -3478
rect 221 -3502 223 -3478
rect 461 -3467 463 -3455
rect 610 -3467 612 -3442
rect 618 -3467 620 -3442
rect 648 -3467 650 -3442
rect 692 -3467 694 -3442
rect 737 -3467 739 -3442
rect 117 -3535 119 -3523
rect 127 -3535 129 -3523
rect 252 -3503 254 -3491
rect 157 -3536 159 -3524
rect 117 -3617 119 -3605
rect 127 -3617 129 -3605
rect 157 -3618 159 -3606
<< ndiffusion >>
rect -76 -2366 -75 -2356
rect -73 -2366 -72 -2356
rect -40 -2366 -39 -2356
rect -37 -2366 -36 -2356
rect -32 -2366 -31 -2356
rect -29 -2366 -28 -2356
rect 4 -2366 5 -2356
rect 7 -2366 8 -2356
rect 12 -2366 13 -2356
rect 15 -2366 16 -2356
rect 55 -2366 56 -2356
rect 58 -2366 59 -2356
rect 529 -2408 530 -2388
rect 532 -2408 533 -2388
rect 235 -2462 236 -2456
rect 238 -2462 239 -2456
rect 492 -2460 493 -2440
rect 495 -2460 496 -2440
rect 194 -2468 195 -2462
rect 197 -2468 199 -2462
rect 203 -2468 205 -2462
rect 207 -2468 208 -2462
rect 562 -2455 563 -2435
rect 565 -2455 566 -2435
rect 830 -2424 831 -2414
rect 833 -2424 834 -2414
rect 866 -2424 867 -2414
rect 869 -2424 870 -2414
rect 874 -2424 875 -2414
rect 877 -2424 878 -2414
rect 910 -2424 911 -2414
rect 913 -2424 914 -2414
rect 918 -2424 919 -2414
rect 921 -2424 922 -2414
rect 961 -2424 962 -2414
rect 964 -2424 965 -2414
rect 605 -2461 606 -2441
rect 608 -2461 609 -2441
rect 95 -2514 96 -2502
rect 98 -2514 106 -2502
rect 108 -2514 109 -2502
rect 135 -2503 136 -2497
rect 138 -2503 139 -2497
rect -839 -2575 -838 -2565
rect -836 -2575 -835 -2565
rect -803 -2575 -802 -2565
rect -800 -2575 -799 -2565
rect -795 -2575 -794 -2565
rect -792 -2575 -791 -2565
rect -759 -2575 -758 -2565
rect -756 -2575 -755 -2565
rect -751 -2575 -750 -2565
rect -748 -2575 -747 -2565
rect -708 -2575 -707 -2565
rect -705 -2575 -704 -2565
rect -626 -2575 -625 -2565
rect -623 -2575 -622 -2565
rect -590 -2575 -589 -2565
rect -587 -2575 -586 -2565
rect -582 -2575 -581 -2565
rect -579 -2575 -578 -2565
rect -546 -2575 -545 -2565
rect -543 -2575 -542 -2565
rect -538 -2575 -537 -2565
rect -535 -2575 -534 -2565
rect -495 -2575 -494 -2565
rect -492 -2575 -491 -2565
rect -338 -2577 -337 -2557
rect -335 -2577 -334 -2557
rect -129 -2582 -128 -2570
rect -126 -2582 -118 -2570
rect -116 -2582 -115 -2570
rect -89 -2571 -88 -2565
rect -86 -2571 -85 -2565
rect -375 -2629 -374 -2609
rect -372 -2629 -371 -2609
rect -305 -2624 -304 -2604
rect -302 -2624 -301 -2604
rect -262 -2630 -261 -2610
rect -259 -2630 -258 -2610
rect 519 -2716 520 -2696
rect 522 -2716 523 -2696
rect 102 -2757 103 -2745
rect 105 -2757 113 -2745
rect 115 -2757 116 -2745
rect 142 -2746 143 -2740
rect 145 -2746 146 -2740
rect 482 -2768 483 -2748
rect 485 -2768 486 -2748
rect 552 -2763 553 -2743
rect 555 -2763 556 -2743
rect 820 -2732 821 -2722
rect 823 -2732 824 -2722
rect 856 -2732 857 -2722
rect 859 -2732 860 -2722
rect 864 -2732 865 -2722
rect 867 -2732 868 -2722
rect 900 -2732 901 -2722
rect 903 -2732 904 -2722
rect 908 -2732 909 -2722
rect 911 -2732 912 -2722
rect 951 -2732 952 -2722
rect 954 -2732 955 -2722
rect 595 -2769 596 -2749
rect 598 -2769 599 -2749
rect 396 -2798 397 -2792
rect 399 -2798 400 -2792
rect 355 -2804 356 -2798
rect 358 -2804 360 -2798
rect 364 -2804 366 -2798
rect 368 -2804 369 -2798
rect 245 -2827 246 -2821
rect 248 -2827 249 -2821
rect 204 -2833 205 -2827
rect 207 -2833 209 -2827
rect 213 -2833 215 -2827
rect 217 -2833 218 -2827
rect -824 -2904 -823 -2894
rect -821 -2904 -820 -2894
rect -788 -2904 -787 -2894
rect -785 -2904 -784 -2894
rect -780 -2904 -779 -2894
rect -777 -2904 -776 -2894
rect -744 -2904 -743 -2894
rect -741 -2904 -740 -2894
rect -736 -2904 -735 -2894
rect -733 -2904 -732 -2894
rect -693 -2904 -692 -2894
rect -690 -2904 -689 -2894
rect -611 -2904 -610 -2894
rect -608 -2904 -607 -2894
rect -575 -2904 -574 -2894
rect -572 -2904 -571 -2894
rect -567 -2904 -566 -2894
rect -564 -2904 -563 -2894
rect -531 -2904 -530 -2894
rect -528 -2904 -527 -2894
rect -523 -2904 -522 -2894
rect -520 -2904 -519 -2894
rect -480 -2904 -479 -2894
rect -477 -2904 -476 -2894
rect -323 -2906 -322 -2886
rect -320 -2906 -319 -2886
rect 105 -2879 106 -2867
rect 108 -2879 116 -2867
rect 118 -2879 119 -2867
rect 145 -2868 146 -2862
rect 148 -2868 149 -2862
rect -114 -2911 -113 -2899
rect -111 -2911 -103 -2899
rect -101 -2911 -100 -2899
rect -74 -2900 -73 -2894
rect -71 -2900 -70 -2894
rect -360 -2958 -359 -2938
rect -357 -2958 -356 -2938
rect -290 -2953 -289 -2933
rect -287 -2953 -286 -2933
rect -247 -2959 -246 -2939
rect -244 -2959 -243 -2939
rect 543 -2975 544 -2955
rect 546 -2975 547 -2955
rect 100 -3021 101 -3009
rect 103 -3021 111 -3009
rect 113 -3021 114 -3009
rect 140 -3010 141 -3004
rect 143 -3010 144 -3004
rect 506 -3027 507 -3007
rect 509 -3027 510 -3007
rect 576 -3022 577 -3002
rect 579 -3022 580 -3002
rect 844 -2991 845 -2981
rect 847 -2991 848 -2981
rect 880 -2991 881 -2981
rect 883 -2991 884 -2981
rect 888 -2991 889 -2981
rect 891 -2991 892 -2981
rect 924 -2991 925 -2981
rect 927 -2991 928 -2981
rect 932 -2991 933 -2981
rect 935 -2991 936 -2981
rect 975 -2991 976 -2981
rect 978 -2991 979 -2981
rect 619 -3028 620 -3008
rect 622 -3028 623 -3008
rect 243 -3091 244 -3085
rect 246 -3091 247 -3085
rect 202 -3097 203 -3091
rect 205 -3097 207 -3091
rect 211 -3097 213 -3091
rect 215 -3097 216 -3091
rect 352 -3118 353 -3112
rect 355 -3118 356 -3112
rect 311 -3124 312 -3118
rect 314 -3124 316 -3118
rect 320 -3124 322 -3118
rect 324 -3124 325 -3118
rect -800 -3171 -799 -3161
rect -797 -3171 -796 -3161
rect -764 -3171 -763 -3161
rect -761 -3171 -760 -3161
rect -756 -3171 -755 -3161
rect -753 -3171 -752 -3161
rect -720 -3171 -719 -3161
rect -717 -3171 -716 -3161
rect -712 -3171 -711 -3161
rect -709 -3171 -708 -3161
rect -669 -3171 -668 -3161
rect -666 -3171 -665 -3161
rect -587 -3171 -586 -3161
rect -584 -3171 -583 -3161
rect -551 -3171 -550 -3161
rect -548 -3171 -547 -3161
rect -543 -3171 -542 -3161
rect -540 -3171 -539 -3161
rect -507 -3171 -506 -3161
rect -504 -3171 -503 -3161
rect -499 -3171 -498 -3161
rect -496 -3171 -495 -3161
rect -456 -3171 -455 -3161
rect -453 -3171 -452 -3161
rect -299 -3173 -298 -3153
rect -296 -3173 -295 -3153
rect 103 -3143 104 -3131
rect 106 -3143 114 -3131
rect 116 -3143 117 -3131
rect 143 -3132 144 -3126
rect 146 -3132 147 -3126
rect -90 -3178 -89 -3166
rect -87 -3178 -79 -3166
rect -77 -3178 -76 -3166
rect -50 -3167 -49 -3161
rect -47 -3167 -46 -3161
rect -336 -3225 -335 -3205
rect -333 -3225 -332 -3205
rect -266 -3220 -265 -3200
rect -263 -3220 -262 -3200
rect 245 -3178 246 -3172
rect 248 -3178 249 -3172
rect -223 -3226 -222 -3206
rect -220 -3226 -219 -3206
rect 204 -3184 205 -3178
rect 207 -3184 209 -3178
rect 213 -3184 215 -3178
rect 217 -3184 218 -3178
rect 110 -3222 111 -3210
rect 113 -3222 121 -3210
rect 123 -3222 124 -3210
rect 150 -3211 151 -3205
rect 153 -3211 154 -3205
rect 564 -3281 565 -3261
rect 567 -3281 568 -3261
rect 527 -3333 528 -3313
rect 530 -3333 531 -3313
rect 597 -3328 598 -3308
rect 600 -3328 601 -3308
rect 865 -3297 866 -3287
rect 868 -3297 869 -3287
rect 901 -3297 902 -3287
rect 904 -3297 905 -3287
rect 909 -3297 910 -3287
rect 912 -3297 913 -3287
rect 945 -3297 946 -3287
rect 948 -3297 949 -3287
rect 953 -3297 954 -3287
rect 956 -3297 957 -3287
rect 996 -3297 997 -3287
rect 999 -3297 1000 -3287
rect 640 -3334 641 -3314
rect 643 -3334 644 -3314
rect 106 -3366 107 -3354
rect 109 -3366 117 -3354
rect 119 -3366 120 -3354
rect 146 -3355 147 -3349
rect 149 -3355 150 -3349
rect 249 -3436 250 -3430
rect 252 -3436 253 -3430
rect -771 -3481 -770 -3471
rect -768 -3481 -767 -3471
rect -735 -3481 -734 -3471
rect -732 -3481 -731 -3471
rect -727 -3481 -726 -3471
rect -724 -3481 -723 -3471
rect -691 -3481 -690 -3471
rect -688 -3481 -687 -3471
rect -683 -3481 -682 -3471
rect -680 -3481 -679 -3471
rect -640 -3481 -639 -3471
rect -637 -3481 -636 -3471
rect -558 -3481 -557 -3471
rect -555 -3481 -554 -3471
rect -522 -3481 -521 -3471
rect -519 -3481 -518 -3471
rect -514 -3481 -513 -3471
rect -511 -3481 -510 -3471
rect -478 -3481 -477 -3471
rect -475 -3481 -474 -3471
rect -470 -3481 -469 -3471
rect -467 -3481 -466 -3471
rect -427 -3481 -426 -3471
rect -424 -3481 -423 -3471
rect 208 -3442 209 -3436
rect 211 -3442 213 -3436
rect 217 -3442 219 -3436
rect 221 -3442 222 -3436
rect -270 -3483 -269 -3463
rect -267 -3483 -266 -3463
rect -61 -3488 -60 -3476
rect -58 -3488 -50 -3476
rect -48 -3488 -47 -3476
rect -21 -3477 -20 -3471
rect -18 -3477 -17 -3471
rect 358 -3463 359 -3457
rect 361 -3463 362 -3457
rect 317 -3469 318 -3463
rect 320 -3469 322 -3463
rect 326 -3469 328 -3463
rect 330 -3469 331 -3463
rect 109 -3488 110 -3476
rect 112 -3488 120 -3476
rect 122 -3488 123 -3476
rect 149 -3477 150 -3471
rect 152 -3477 153 -3471
rect -307 -3535 -306 -3515
rect -304 -3535 -303 -3515
rect -237 -3530 -236 -3510
rect -234 -3530 -233 -3510
rect 460 -3487 461 -3481
rect 463 -3487 464 -3481
rect -194 -3536 -193 -3516
rect -191 -3536 -190 -3516
rect 419 -3493 420 -3487
rect 422 -3493 424 -3487
rect 428 -3493 430 -3487
rect 432 -3493 433 -3487
rect 605 -3499 606 -3489
rect 608 -3499 609 -3489
rect 641 -3499 642 -3489
rect 644 -3499 645 -3489
rect 649 -3499 650 -3489
rect 652 -3499 653 -3489
rect 685 -3499 686 -3489
rect 688 -3499 689 -3489
rect 693 -3499 694 -3489
rect 696 -3499 697 -3489
rect 736 -3499 737 -3489
rect 739 -3499 740 -3489
rect 251 -3523 252 -3517
rect 254 -3523 255 -3517
rect 210 -3529 211 -3523
rect 213 -3529 215 -3523
rect 219 -3529 221 -3523
rect 223 -3529 224 -3523
rect 116 -3567 117 -3555
rect 119 -3567 127 -3555
rect 129 -3567 130 -3555
rect 156 -3556 157 -3550
rect 159 -3556 160 -3550
rect 116 -3649 117 -3637
rect 119 -3649 127 -3637
rect 129 -3649 130 -3637
rect 156 -3638 157 -3632
rect 159 -3638 160 -3632
<< pdiffusion >>
rect -72 -2334 -71 -2309
rect -69 -2334 -68 -2309
rect -64 -2334 -63 -2309
rect -61 -2334 -60 -2309
rect -34 -2334 -33 -2309
rect -31 -2334 -30 -2309
rect 10 -2334 11 -2309
rect 13 -2334 14 -2309
rect 55 -2334 56 -2309
rect 58 -2334 59 -2309
rect 194 -2441 195 -2417
rect 197 -2441 205 -2417
rect 207 -2441 208 -2417
rect 492 -2420 493 -2380
rect 495 -2420 496 -2380
rect 562 -2415 563 -2395
rect 565 -2415 566 -2395
rect 235 -2442 236 -2430
rect 238 -2442 239 -2430
rect 605 -2421 606 -2381
rect 608 -2421 609 -2381
rect 834 -2392 835 -2367
rect 837 -2392 838 -2367
rect 842 -2392 843 -2367
rect 845 -2392 846 -2367
rect 872 -2392 873 -2367
rect 875 -2392 876 -2367
rect 916 -2392 917 -2367
rect 919 -2392 920 -2367
rect 961 -2392 962 -2367
rect 964 -2392 965 -2367
rect 529 -2448 530 -2428
rect 532 -2448 533 -2428
rect 95 -2482 96 -2470
rect 98 -2482 100 -2470
rect 104 -2482 106 -2470
rect 108 -2482 109 -2470
rect 135 -2483 136 -2471
rect 138 -2483 139 -2471
rect -835 -2543 -834 -2518
rect -832 -2543 -831 -2518
rect -827 -2543 -826 -2518
rect -824 -2543 -823 -2518
rect -797 -2543 -796 -2518
rect -794 -2543 -793 -2518
rect -753 -2543 -752 -2518
rect -750 -2543 -749 -2518
rect -708 -2543 -707 -2518
rect -705 -2543 -704 -2518
rect -622 -2543 -621 -2518
rect -619 -2543 -618 -2518
rect -614 -2543 -613 -2518
rect -611 -2543 -610 -2518
rect -584 -2543 -583 -2518
rect -581 -2543 -580 -2518
rect -540 -2543 -539 -2518
rect -537 -2543 -536 -2518
rect -495 -2543 -494 -2518
rect -492 -2543 -491 -2518
rect -375 -2589 -374 -2549
rect -372 -2589 -371 -2549
rect -129 -2550 -128 -2538
rect -126 -2550 -124 -2538
rect -120 -2550 -118 -2538
rect -116 -2550 -115 -2538
rect -305 -2584 -304 -2564
rect -302 -2584 -301 -2564
rect -262 -2590 -261 -2550
rect -259 -2590 -258 -2550
rect -89 -2551 -88 -2539
rect -86 -2551 -85 -2539
rect -338 -2617 -337 -2597
rect -335 -2617 -334 -2597
rect 102 -2725 103 -2713
rect 105 -2725 107 -2713
rect 111 -2725 113 -2713
rect 115 -2725 116 -2713
rect 142 -2726 143 -2714
rect 145 -2726 146 -2714
rect 482 -2728 483 -2688
rect 485 -2728 486 -2688
rect 552 -2723 553 -2703
rect 555 -2723 556 -2703
rect 595 -2729 596 -2689
rect 598 -2729 599 -2689
rect 824 -2700 825 -2675
rect 827 -2700 828 -2675
rect 832 -2700 833 -2675
rect 835 -2700 836 -2675
rect 862 -2700 863 -2675
rect 865 -2700 866 -2675
rect 906 -2700 907 -2675
rect 909 -2700 910 -2675
rect 951 -2700 952 -2675
rect 954 -2700 955 -2675
rect 355 -2777 356 -2753
rect 358 -2777 366 -2753
rect 368 -2777 369 -2753
rect 204 -2806 205 -2782
rect 207 -2806 215 -2782
rect 217 -2806 218 -2782
rect 245 -2807 246 -2795
rect 248 -2807 249 -2795
rect 396 -2778 397 -2766
rect 399 -2778 400 -2766
rect 519 -2756 520 -2736
rect 522 -2756 523 -2736
rect 105 -2847 106 -2835
rect 108 -2847 110 -2835
rect 114 -2847 116 -2835
rect 118 -2847 119 -2835
rect -820 -2872 -819 -2847
rect -817 -2872 -816 -2847
rect -812 -2872 -811 -2847
rect -809 -2872 -808 -2847
rect -782 -2872 -781 -2847
rect -779 -2872 -778 -2847
rect -738 -2872 -737 -2847
rect -735 -2872 -734 -2847
rect -693 -2872 -692 -2847
rect -690 -2872 -689 -2847
rect -607 -2872 -606 -2847
rect -604 -2872 -603 -2847
rect -599 -2872 -598 -2847
rect -596 -2872 -595 -2847
rect -569 -2872 -568 -2847
rect -566 -2872 -565 -2847
rect -525 -2872 -524 -2847
rect -522 -2872 -521 -2847
rect -480 -2872 -479 -2847
rect -477 -2872 -476 -2847
rect -360 -2918 -359 -2878
rect -357 -2918 -356 -2878
rect -114 -2879 -113 -2867
rect -111 -2879 -109 -2867
rect -105 -2879 -103 -2867
rect -101 -2879 -100 -2867
rect 145 -2848 146 -2836
rect 148 -2848 149 -2836
rect -290 -2913 -289 -2893
rect -287 -2913 -286 -2893
rect -247 -2919 -246 -2879
rect -244 -2919 -243 -2879
rect -74 -2880 -73 -2868
rect -71 -2880 -70 -2868
rect -323 -2946 -322 -2926
rect -320 -2946 -319 -2926
rect 100 -2989 101 -2977
rect 103 -2989 105 -2977
rect 109 -2989 111 -2977
rect 113 -2989 114 -2977
rect 140 -2990 141 -2978
rect 143 -2990 144 -2978
rect 506 -2987 507 -2947
rect 509 -2987 510 -2947
rect 576 -2982 577 -2962
rect 579 -2982 580 -2962
rect 619 -2988 620 -2948
rect 622 -2988 623 -2948
rect 848 -2959 849 -2934
rect 851 -2959 852 -2934
rect 856 -2959 857 -2934
rect 859 -2959 860 -2934
rect 886 -2959 887 -2934
rect 889 -2959 890 -2934
rect 930 -2959 931 -2934
rect 933 -2959 934 -2934
rect 975 -2959 976 -2934
rect 978 -2959 979 -2934
rect 543 -3015 544 -2995
rect 546 -3015 547 -2995
rect 202 -3070 203 -3046
rect 205 -3070 213 -3046
rect 215 -3070 216 -3046
rect 243 -3071 244 -3059
rect 246 -3071 247 -3059
rect 311 -3097 312 -3073
rect 314 -3097 322 -3073
rect 324 -3097 325 -3073
rect 103 -3111 104 -3099
rect 106 -3111 108 -3099
rect 112 -3111 114 -3099
rect 116 -3111 117 -3099
rect -796 -3139 -795 -3114
rect -793 -3139 -792 -3114
rect -788 -3139 -787 -3114
rect -785 -3139 -784 -3114
rect -758 -3139 -757 -3114
rect -755 -3139 -754 -3114
rect -714 -3139 -713 -3114
rect -711 -3139 -710 -3114
rect -669 -3139 -668 -3114
rect -666 -3139 -665 -3114
rect -583 -3139 -582 -3114
rect -580 -3139 -579 -3114
rect -575 -3139 -574 -3114
rect -572 -3139 -571 -3114
rect -545 -3139 -544 -3114
rect -542 -3139 -541 -3114
rect -501 -3139 -500 -3114
rect -498 -3139 -497 -3114
rect -456 -3139 -455 -3114
rect -453 -3139 -452 -3114
rect 143 -3112 144 -3100
rect 146 -3112 147 -3100
rect 352 -3098 353 -3086
rect 355 -3098 356 -3086
rect -336 -3185 -335 -3145
rect -333 -3185 -332 -3145
rect -90 -3146 -89 -3134
rect -87 -3146 -85 -3134
rect -81 -3146 -79 -3134
rect -77 -3146 -76 -3134
rect -266 -3180 -265 -3160
rect -263 -3180 -262 -3160
rect -223 -3186 -222 -3146
rect -220 -3186 -219 -3146
rect -50 -3147 -49 -3135
rect -47 -3147 -46 -3135
rect 204 -3157 205 -3133
rect 207 -3157 215 -3133
rect 217 -3157 218 -3133
rect -299 -3213 -298 -3193
rect -296 -3213 -295 -3193
rect 110 -3190 111 -3178
rect 113 -3190 115 -3178
rect 119 -3190 121 -3178
rect 123 -3190 124 -3178
rect 245 -3158 246 -3146
rect 248 -3158 249 -3146
rect 150 -3191 151 -3179
rect 153 -3191 154 -3179
rect 527 -3293 528 -3253
rect 530 -3293 531 -3253
rect 597 -3288 598 -3268
rect 600 -3288 601 -3268
rect 640 -3294 641 -3254
rect 643 -3294 644 -3254
rect 869 -3265 870 -3240
rect 872 -3265 873 -3240
rect 877 -3265 878 -3240
rect 880 -3265 881 -3240
rect 907 -3265 908 -3240
rect 910 -3265 911 -3240
rect 951 -3265 952 -3240
rect 954 -3265 955 -3240
rect 996 -3265 997 -3240
rect 999 -3265 1000 -3240
rect 106 -3334 107 -3322
rect 109 -3334 111 -3322
rect 115 -3334 117 -3322
rect 119 -3334 120 -3322
rect 146 -3335 147 -3323
rect 149 -3335 150 -3323
rect 564 -3321 565 -3301
rect 567 -3321 568 -3301
rect 208 -3415 209 -3391
rect 211 -3415 219 -3391
rect 221 -3415 222 -3391
rect -767 -3449 -766 -3424
rect -764 -3449 -763 -3424
rect -759 -3449 -758 -3424
rect -756 -3449 -755 -3424
rect -729 -3449 -728 -3424
rect -726 -3449 -725 -3424
rect -685 -3449 -684 -3424
rect -682 -3449 -681 -3424
rect -640 -3449 -639 -3424
rect -637 -3449 -636 -3424
rect -554 -3449 -553 -3424
rect -551 -3449 -550 -3424
rect -546 -3449 -545 -3424
rect -543 -3449 -542 -3424
rect -516 -3449 -515 -3424
rect -513 -3449 -512 -3424
rect -472 -3449 -471 -3424
rect -469 -3449 -468 -3424
rect -427 -3449 -426 -3424
rect -424 -3449 -423 -3424
rect 249 -3416 250 -3404
rect 252 -3416 253 -3404
rect -307 -3495 -306 -3455
rect -304 -3495 -303 -3455
rect -61 -3456 -60 -3444
rect -58 -3456 -56 -3444
rect -52 -3456 -50 -3444
rect -48 -3456 -47 -3444
rect 317 -3442 318 -3418
rect 320 -3442 328 -3418
rect 330 -3442 331 -3418
rect -237 -3490 -236 -3470
rect -234 -3490 -233 -3470
rect -194 -3496 -193 -3456
rect -191 -3496 -190 -3456
rect -21 -3457 -20 -3445
rect -18 -3457 -17 -3445
rect 109 -3456 110 -3444
rect 112 -3456 114 -3444
rect 118 -3456 120 -3444
rect 122 -3456 123 -3444
rect 149 -3457 150 -3445
rect 152 -3457 153 -3445
rect 358 -3443 359 -3431
rect 361 -3443 362 -3431
rect 419 -3466 420 -3442
rect 422 -3466 430 -3442
rect 432 -3466 433 -3442
rect -270 -3523 -269 -3503
rect -267 -3523 -266 -3503
rect 210 -3502 211 -3478
rect 213 -3502 221 -3478
rect 223 -3502 224 -3478
rect 460 -3467 461 -3455
rect 463 -3467 464 -3455
rect 609 -3467 610 -3442
rect 612 -3467 613 -3442
rect 617 -3467 618 -3442
rect 620 -3467 621 -3442
rect 647 -3467 648 -3442
rect 650 -3467 651 -3442
rect 691 -3467 692 -3442
rect 694 -3467 695 -3442
rect 736 -3467 737 -3442
rect 739 -3467 740 -3442
rect 116 -3535 117 -3523
rect 119 -3535 121 -3523
rect 125 -3535 127 -3523
rect 129 -3535 130 -3523
rect 251 -3503 252 -3491
rect 254 -3503 255 -3491
rect 156 -3536 157 -3524
rect 159 -3536 160 -3524
rect 116 -3617 117 -3605
rect 119 -3617 121 -3605
rect 125 -3617 127 -3605
rect 129 -3617 130 -3605
rect 156 -3618 157 -3606
rect 159 -3618 160 -3606
<< ndcontact >>
rect -80 -2366 -76 -2356
rect -72 -2366 -68 -2356
rect -44 -2366 -40 -2356
rect -36 -2366 -32 -2356
rect -28 -2366 -24 -2356
rect 0 -2366 4 -2356
rect 8 -2366 12 -2356
rect 16 -2366 20 -2356
rect 51 -2366 55 -2356
rect 59 -2366 63 -2356
rect 525 -2408 529 -2388
rect 533 -2408 537 -2388
rect 231 -2462 235 -2456
rect 239 -2462 243 -2456
rect 488 -2460 492 -2440
rect 496 -2460 500 -2440
rect 190 -2468 194 -2462
rect 199 -2468 203 -2462
rect 208 -2468 212 -2462
rect 558 -2455 562 -2435
rect 566 -2455 570 -2435
rect 826 -2424 830 -2414
rect 834 -2424 838 -2414
rect 862 -2424 866 -2414
rect 870 -2424 874 -2414
rect 878 -2424 882 -2414
rect 906 -2424 910 -2414
rect 914 -2424 918 -2414
rect 922 -2424 926 -2414
rect 957 -2424 961 -2414
rect 965 -2424 969 -2414
rect 601 -2461 605 -2441
rect 609 -2461 613 -2441
rect 91 -2514 95 -2502
rect 109 -2514 113 -2502
rect 131 -2503 135 -2497
rect 139 -2503 143 -2497
rect -843 -2575 -839 -2565
rect -835 -2575 -831 -2565
rect -807 -2575 -803 -2565
rect -799 -2575 -795 -2565
rect -791 -2575 -787 -2565
rect -763 -2575 -759 -2565
rect -755 -2575 -751 -2565
rect -747 -2575 -743 -2565
rect -712 -2575 -708 -2565
rect -704 -2575 -700 -2565
rect -630 -2575 -626 -2565
rect -622 -2575 -618 -2565
rect -594 -2575 -590 -2565
rect -586 -2575 -582 -2565
rect -578 -2575 -574 -2565
rect -550 -2575 -546 -2565
rect -542 -2575 -538 -2565
rect -534 -2575 -530 -2565
rect -499 -2575 -495 -2565
rect -491 -2575 -487 -2565
rect -342 -2577 -338 -2557
rect -334 -2577 -330 -2557
rect -133 -2582 -129 -2570
rect -115 -2582 -111 -2570
rect -93 -2571 -89 -2565
rect -85 -2571 -81 -2565
rect -379 -2629 -375 -2609
rect -371 -2629 -367 -2609
rect -309 -2624 -305 -2604
rect -301 -2624 -297 -2604
rect -266 -2630 -262 -2610
rect -258 -2630 -254 -2610
rect 515 -2716 519 -2696
rect 523 -2716 527 -2696
rect 98 -2757 102 -2745
rect 116 -2757 120 -2745
rect 138 -2746 142 -2740
rect 146 -2746 150 -2740
rect 478 -2768 482 -2748
rect 486 -2768 490 -2748
rect 548 -2763 552 -2743
rect 556 -2763 560 -2743
rect 816 -2732 820 -2722
rect 824 -2732 828 -2722
rect 852 -2732 856 -2722
rect 860 -2732 864 -2722
rect 868 -2732 872 -2722
rect 896 -2732 900 -2722
rect 904 -2732 908 -2722
rect 912 -2732 916 -2722
rect 947 -2732 951 -2722
rect 955 -2732 959 -2722
rect 591 -2769 595 -2749
rect 599 -2769 603 -2749
rect 392 -2798 396 -2792
rect 400 -2798 404 -2792
rect 351 -2804 355 -2798
rect 360 -2804 364 -2798
rect 369 -2804 373 -2798
rect 241 -2827 245 -2821
rect 249 -2827 253 -2821
rect 200 -2833 204 -2827
rect 209 -2833 213 -2827
rect 218 -2833 222 -2827
rect -828 -2904 -824 -2894
rect -820 -2904 -816 -2894
rect -792 -2904 -788 -2894
rect -784 -2904 -780 -2894
rect -776 -2904 -772 -2894
rect -748 -2904 -744 -2894
rect -740 -2904 -736 -2894
rect -732 -2904 -728 -2894
rect -697 -2904 -693 -2894
rect -689 -2904 -685 -2894
rect -615 -2904 -611 -2894
rect -607 -2904 -603 -2894
rect -579 -2904 -575 -2894
rect -571 -2904 -567 -2894
rect -563 -2904 -559 -2894
rect -535 -2904 -531 -2894
rect -527 -2904 -523 -2894
rect -519 -2904 -515 -2894
rect -484 -2904 -480 -2894
rect -476 -2904 -472 -2894
rect -327 -2906 -323 -2886
rect -319 -2906 -315 -2886
rect 101 -2879 105 -2867
rect 119 -2879 123 -2867
rect 141 -2868 145 -2862
rect 149 -2868 153 -2862
rect -118 -2911 -114 -2899
rect -100 -2911 -96 -2899
rect -78 -2900 -74 -2894
rect -70 -2900 -66 -2894
rect -364 -2958 -360 -2938
rect -356 -2958 -352 -2938
rect -294 -2953 -290 -2933
rect -286 -2953 -282 -2933
rect -251 -2959 -247 -2939
rect -243 -2959 -239 -2939
rect 539 -2975 543 -2955
rect 547 -2975 551 -2955
rect 96 -3021 100 -3009
rect 114 -3021 118 -3009
rect 136 -3010 140 -3004
rect 144 -3010 148 -3004
rect 502 -3027 506 -3007
rect 510 -3027 514 -3007
rect 572 -3022 576 -3002
rect 580 -3022 584 -3002
rect 840 -2991 844 -2981
rect 848 -2991 852 -2981
rect 876 -2991 880 -2981
rect 884 -2991 888 -2981
rect 892 -2991 896 -2981
rect 920 -2991 924 -2981
rect 928 -2991 932 -2981
rect 936 -2991 940 -2981
rect 971 -2991 975 -2981
rect 979 -2991 983 -2981
rect 615 -3028 619 -3008
rect 623 -3028 627 -3008
rect 239 -3091 243 -3085
rect 247 -3091 251 -3085
rect 198 -3097 202 -3091
rect 207 -3097 211 -3091
rect 216 -3097 220 -3091
rect 348 -3118 352 -3112
rect 356 -3118 360 -3112
rect 307 -3124 311 -3118
rect 316 -3124 320 -3118
rect 325 -3124 329 -3118
rect -804 -3171 -800 -3161
rect -796 -3171 -792 -3161
rect -768 -3171 -764 -3161
rect -760 -3171 -756 -3161
rect -752 -3171 -748 -3161
rect -724 -3171 -720 -3161
rect -716 -3171 -712 -3161
rect -708 -3171 -704 -3161
rect -673 -3171 -669 -3161
rect -665 -3171 -661 -3161
rect -591 -3171 -587 -3161
rect -583 -3171 -579 -3161
rect -555 -3171 -551 -3161
rect -547 -3171 -543 -3161
rect -539 -3171 -535 -3161
rect -511 -3171 -507 -3161
rect -503 -3171 -499 -3161
rect -495 -3171 -491 -3161
rect -460 -3171 -456 -3161
rect -452 -3171 -448 -3161
rect -303 -3173 -299 -3153
rect -295 -3173 -291 -3153
rect 99 -3143 103 -3131
rect 117 -3143 121 -3131
rect 139 -3132 143 -3126
rect 147 -3132 151 -3126
rect -94 -3178 -90 -3166
rect -76 -3178 -72 -3166
rect -54 -3167 -50 -3161
rect -46 -3167 -42 -3161
rect -340 -3225 -336 -3205
rect -332 -3225 -328 -3205
rect -270 -3220 -266 -3200
rect -262 -3220 -258 -3200
rect 241 -3178 245 -3172
rect 249 -3178 253 -3172
rect -227 -3226 -223 -3206
rect -219 -3226 -215 -3206
rect 200 -3184 204 -3178
rect 209 -3184 213 -3178
rect 218 -3184 222 -3178
rect 106 -3222 110 -3210
rect 124 -3222 128 -3210
rect 146 -3211 150 -3205
rect 154 -3211 158 -3205
rect 560 -3281 564 -3261
rect 568 -3281 572 -3261
rect 523 -3333 527 -3313
rect 531 -3333 535 -3313
rect 593 -3328 597 -3308
rect 601 -3328 605 -3308
rect 861 -3297 865 -3287
rect 869 -3297 873 -3287
rect 897 -3297 901 -3287
rect 905 -3297 909 -3287
rect 913 -3297 917 -3287
rect 941 -3297 945 -3287
rect 949 -3297 953 -3287
rect 957 -3297 961 -3287
rect 992 -3297 996 -3287
rect 1000 -3297 1004 -3287
rect 636 -3334 640 -3314
rect 644 -3334 648 -3314
rect 102 -3366 106 -3354
rect 120 -3366 124 -3354
rect 142 -3355 146 -3349
rect 150 -3355 154 -3349
rect 245 -3436 249 -3430
rect 253 -3436 257 -3430
rect -775 -3481 -771 -3471
rect -767 -3481 -763 -3471
rect -739 -3481 -735 -3471
rect -731 -3481 -727 -3471
rect -723 -3481 -719 -3471
rect -695 -3481 -691 -3471
rect -687 -3481 -683 -3471
rect -679 -3481 -675 -3471
rect -644 -3481 -640 -3471
rect -636 -3481 -632 -3471
rect -562 -3481 -558 -3471
rect -554 -3481 -550 -3471
rect -526 -3481 -522 -3471
rect -518 -3481 -514 -3471
rect -510 -3481 -506 -3471
rect -482 -3481 -478 -3471
rect -474 -3481 -470 -3471
rect -466 -3481 -462 -3471
rect -431 -3481 -427 -3471
rect -423 -3481 -419 -3471
rect 204 -3442 208 -3436
rect 213 -3442 217 -3436
rect 222 -3442 226 -3436
rect -274 -3483 -270 -3463
rect -266 -3483 -262 -3463
rect -65 -3488 -61 -3476
rect -47 -3488 -43 -3476
rect -25 -3477 -21 -3471
rect -17 -3477 -13 -3471
rect 354 -3463 358 -3457
rect 362 -3463 366 -3457
rect 313 -3469 317 -3463
rect 322 -3469 326 -3463
rect 331 -3469 335 -3463
rect 105 -3488 109 -3476
rect 123 -3488 127 -3476
rect 145 -3477 149 -3471
rect 153 -3477 157 -3471
rect -311 -3535 -307 -3515
rect -303 -3535 -299 -3515
rect -241 -3530 -237 -3510
rect -233 -3530 -229 -3510
rect 456 -3487 460 -3481
rect 464 -3487 468 -3481
rect -198 -3536 -194 -3516
rect -190 -3536 -186 -3516
rect 415 -3493 419 -3487
rect 424 -3493 428 -3487
rect 433 -3493 437 -3487
rect 601 -3499 605 -3489
rect 609 -3499 613 -3489
rect 637 -3499 641 -3489
rect 645 -3499 649 -3489
rect 653 -3499 657 -3489
rect 681 -3499 685 -3489
rect 689 -3499 693 -3489
rect 697 -3499 701 -3489
rect 732 -3499 736 -3489
rect 740 -3499 744 -3489
rect 247 -3523 251 -3517
rect 255 -3523 259 -3517
rect 206 -3529 210 -3523
rect 215 -3529 219 -3523
rect 224 -3529 228 -3523
rect 112 -3567 116 -3555
rect 130 -3567 134 -3555
rect 152 -3556 156 -3550
rect 160 -3556 164 -3550
rect 112 -3649 116 -3637
rect 130 -3649 134 -3637
rect 152 -3638 156 -3632
rect 160 -3638 164 -3632
<< pdcontact >>
rect -76 -2334 -72 -2309
rect -68 -2334 -64 -2309
rect -60 -2334 -56 -2309
rect -38 -2334 -34 -2309
rect -30 -2334 -26 -2309
rect 6 -2334 10 -2309
rect 14 -2334 18 -2309
rect 51 -2334 55 -2309
rect 59 -2334 63 -2309
rect 190 -2441 194 -2417
rect 208 -2441 212 -2417
rect 488 -2420 492 -2380
rect 496 -2420 500 -2380
rect 558 -2415 562 -2395
rect 566 -2415 570 -2395
rect 231 -2442 235 -2430
rect 239 -2442 243 -2430
rect 601 -2421 605 -2381
rect 609 -2421 613 -2381
rect 830 -2392 834 -2367
rect 838 -2392 842 -2367
rect 846 -2392 850 -2367
rect 868 -2392 872 -2367
rect 876 -2392 880 -2367
rect 912 -2392 916 -2367
rect 920 -2392 924 -2367
rect 957 -2392 961 -2367
rect 965 -2392 969 -2367
rect 525 -2448 529 -2428
rect 533 -2448 537 -2428
rect 91 -2482 95 -2470
rect 100 -2482 104 -2470
rect 109 -2482 113 -2470
rect 131 -2483 135 -2471
rect 139 -2483 143 -2471
rect -839 -2543 -835 -2518
rect -831 -2543 -827 -2518
rect -823 -2543 -819 -2518
rect -801 -2543 -797 -2518
rect -793 -2543 -789 -2518
rect -757 -2543 -753 -2518
rect -749 -2543 -745 -2518
rect -712 -2543 -708 -2518
rect -704 -2543 -700 -2518
rect -626 -2543 -622 -2518
rect -618 -2543 -614 -2518
rect -610 -2543 -606 -2518
rect -588 -2543 -584 -2518
rect -580 -2543 -576 -2518
rect -544 -2543 -540 -2518
rect -536 -2543 -532 -2518
rect -499 -2543 -495 -2518
rect -491 -2543 -487 -2518
rect -379 -2589 -375 -2549
rect -371 -2589 -367 -2549
rect -133 -2550 -129 -2538
rect -124 -2550 -120 -2538
rect -115 -2550 -111 -2538
rect -309 -2584 -305 -2564
rect -301 -2584 -297 -2564
rect -266 -2590 -262 -2550
rect -258 -2590 -254 -2550
rect -93 -2551 -89 -2539
rect -85 -2551 -81 -2539
rect -342 -2617 -338 -2597
rect -334 -2617 -330 -2597
rect 98 -2725 102 -2713
rect 107 -2725 111 -2713
rect 116 -2725 120 -2713
rect 138 -2726 142 -2714
rect 146 -2726 150 -2714
rect 478 -2728 482 -2688
rect 486 -2728 490 -2688
rect 548 -2723 552 -2703
rect 556 -2723 560 -2703
rect 591 -2729 595 -2689
rect 599 -2729 603 -2689
rect 820 -2700 824 -2675
rect 828 -2700 832 -2675
rect 836 -2700 840 -2675
rect 858 -2700 862 -2675
rect 866 -2700 870 -2675
rect 902 -2700 906 -2675
rect 910 -2700 914 -2675
rect 947 -2700 951 -2675
rect 955 -2700 959 -2675
rect 351 -2777 355 -2753
rect 369 -2777 373 -2753
rect 200 -2806 204 -2782
rect 218 -2806 222 -2782
rect 241 -2807 245 -2795
rect 249 -2807 253 -2795
rect 392 -2778 396 -2766
rect 400 -2778 404 -2766
rect 515 -2756 519 -2736
rect 523 -2756 527 -2736
rect 101 -2847 105 -2835
rect 110 -2847 114 -2835
rect 119 -2847 123 -2835
rect -824 -2872 -820 -2847
rect -816 -2872 -812 -2847
rect -808 -2872 -804 -2847
rect -786 -2872 -782 -2847
rect -778 -2872 -774 -2847
rect -742 -2872 -738 -2847
rect -734 -2872 -730 -2847
rect -697 -2872 -693 -2847
rect -689 -2872 -685 -2847
rect -611 -2872 -607 -2847
rect -603 -2872 -599 -2847
rect -595 -2872 -591 -2847
rect -573 -2872 -569 -2847
rect -565 -2872 -561 -2847
rect -529 -2872 -525 -2847
rect -521 -2872 -517 -2847
rect -484 -2872 -480 -2847
rect -476 -2872 -472 -2847
rect -364 -2918 -360 -2878
rect -356 -2918 -352 -2878
rect -118 -2879 -114 -2867
rect -109 -2879 -105 -2867
rect -100 -2879 -96 -2867
rect 141 -2848 145 -2836
rect 149 -2848 153 -2836
rect -294 -2913 -290 -2893
rect -286 -2913 -282 -2893
rect -251 -2919 -247 -2879
rect -243 -2919 -239 -2879
rect -78 -2880 -74 -2868
rect -70 -2880 -66 -2868
rect -327 -2946 -323 -2926
rect -319 -2946 -315 -2926
rect 96 -2989 100 -2977
rect 105 -2989 109 -2977
rect 114 -2989 118 -2977
rect 136 -2990 140 -2978
rect 144 -2990 148 -2978
rect 502 -2987 506 -2947
rect 510 -2987 514 -2947
rect 572 -2982 576 -2962
rect 580 -2982 584 -2962
rect 615 -2988 619 -2948
rect 623 -2988 627 -2948
rect 844 -2959 848 -2934
rect 852 -2959 856 -2934
rect 860 -2959 864 -2934
rect 882 -2959 886 -2934
rect 890 -2959 894 -2934
rect 926 -2959 930 -2934
rect 934 -2959 938 -2934
rect 971 -2959 975 -2934
rect 979 -2959 983 -2934
rect 539 -3015 543 -2995
rect 547 -3015 551 -2995
rect 198 -3070 202 -3046
rect 216 -3070 220 -3046
rect 239 -3071 243 -3059
rect 247 -3071 251 -3059
rect 307 -3097 311 -3073
rect 325 -3097 329 -3073
rect 99 -3111 103 -3099
rect 108 -3111 112 -3099
rect 117 -3111 121 -3099
rect -800 -3139 -796 -3114
rect -792 -3139 -788 -3114
rect -784 -3139 -780 -3114
rect -762 -3139 -758 -3114
rect -754 -3139 -750 -3114
rect -718 -3139 -714 -3114
rect -710 -3139 -706 -3114
rect -673 -3139 -669 -3114
rect -665 -3139 -661 -3114
rect -587 -3139 -583 -3114
rect -579 -3139 -575 -3114
rect -571 -3139 -567 -3114
rect -549 -3139 -545 -3114
rect -541 -3139 -537 -3114
rect -505 -3139 -501 -3114
rect -497 -3139 -493 -3114
rect -460 -3139 -456 -3114
rect -452 -3139 -448 -3114
rect 139 -3112 143 -3100
rect 147 -3112 151 -3100
rect 348 -3098 352 -3086
rect 356 -3098 360 -3086
rect -340 -3185 -336 -3145
rect -332 -3185 -328 -3145
rect -94 -3146 -90 -3134
rect -85 -3146 -81 -3134
rect -76 -3146 -72 -3134
rect -270 -3180 -266 -3160
rect -262 -3180 -258 -3160
rect -227 -3186 -223 -3146
rect -219 -3186 -215 -3146
rect -54 -3147 -50 -3135
rect -46 -3147 -42 -3135
rect 200 -3157 204 -3133
rect 218 -3157 222 -3133
rect -303 -3213 -299 -3193
rect -295 -3213 -291 -3193
rect 106 -3190 110 -3178
rect 115 -3190 119 -3178
rect 124 -3190 128 -3178
rect 241 -3158 245 -3146
rect 249 -3158 253 -3146
rect 146 -3191 150 -3179
rect 154 -3191 158 -3179
rect 523 -3293 527 -3253
rect 531 -3293 535 -3253
rect 593 -3288 597 -3268
rect 601 -3288 605 -3268
rect 636 -3294 640 -3254
rect 644 -3294 648 -3254
rect 865 -3265 869 -3240
rect 873 -3265 877 -3240
rect 881 -3265 885 -3240
rect 903 -3265 907 -3240
rect 911 -3265 915 -3240
rect 947 -3265 951 -3240
rect 955 -3265 959 -3240
rect 992 -3265 996 -3240
rect 1000 -3265 1004 -3240
rect 102 -3334 106 -3322
rect 111 -3334 115 -3322
rect 120 -3334 124 -3322
rect 142 -3335 146 -3323
rect 150 -3335 154 -3323
rect 560 -3321 564 -3301
rect 568 -3321 572 -3301
rect 204 -3415 208 -3391
rect 222 -3415 226 -3391
rect -771 -3449 -767 -3424
rect -763 -3449 -759 -3424
rect -755 -3449 -751 -3424
rect -733 -3449 -729 -3424
rect -725 -3449 -721 -3424
rect -689 -3449 -685 -3424
rect -681 -3449 -677 -3424
rect -644 -3449 -640 -3424
rect -636 -3449 -632 -3424
rect -558 -3449 -554 -3424
rect -550 -3449 -546 -3424
rect -542 -3449 -538 -3424
rect -520 -3449 -516 -3424
rect -512 -3449 -508 -3424
rect -476 -3449 -472 -3424
rect -468 -3449 -464 -3424
rect -431 -3449 -427 -3424
rect -423 -3449 -419 -3424
rect 245 -3416 249 -3404
rect 253 -3416 257 -3404
rect -311 -3495 -307 -3455
rect -303 -3495 -299 -3455
rect -65 -3456 -61 -3444
rect -56 -3456 -52 -3444
rect -47 -3456 -43 -3444
rect 313 -3442 317 -3418
rect 331 -3442 335 -3418
rect -241 -3490 -237 -3470
rect -233 -3490 -229 -3470
rect -198 -3496 -194 -3456
rect -190 -3496 -186 -3456
rect -25 -3457 -21 -3445
rect -17 -3457 -13 -3445
rect 105 -3456 109 -3444
rect 114 -3456 118 -3444
rect 123 -3456 127 -3444
rect 145 -3457 149 -3445
rect 153 -3457 157 -3445
rect 354 -3443 358 -3431
rect 362 -3443 366 -3431
rect 415 -3466 419 -3442
rect 433 -3466 437 -3442
rect -274 -3523 -270 -3503
rect -266 -3523 -262 -3503
rect 206 -3502 210 -3478
rect 224 -3502 228 -3478
rect 456 -3467 460 -3455
rect 464 -3467 468 -3455
rect 605 -3467 609 -3442
rect 613 -3467 617 -3442
rect 621 -3467 625 -3442
rect 643 -3467 647 -3442
rect 651 -3467 655 -3442
rect 687 -3467 691 -3442
rect 695 -3467 699 -3442
rect 732 -3467 736 -3442
rect 740 -3467 744 -3442
rect 112 -3535 116 -3523
rect 121 -3535 125 -3523
rect 130 -3535 134 -3523
rect 247 -3503 251 -3491
rect 255 -3503 259 -3491
rect 152 -3536 156 -3524
rect 160 -3536 164 -3524
rect 112 -3617 116 -3605
rect 121 -3617 125 -3605
rect 130 -3617 134 -3605
rect 152 -3618 156 -3606
rect 160 -3618 164 -3606
<< polysilicon >>
rect -71 -2309 -69 -2306
rect -63 -2309 -61 -2306
rect -33 -2309 -31 -2306
rect 11 -2309 13 -2306
rect 56 -2309 58 -2306
rect -71 -2341 -69 -2334
rect -76 -2345 -69 -2341
rect -75 -2356 -73 -2345
rect -63 -2353 -61 -2334
rect -33 -2342 -31 -2334
rect 11 -2342 13 -2334
rect -39 -2344 -31 -2342
rect 5 -2344 13 -2342
rect -39 -2356 -37 -2344
rect -31 -2356 -29 -2347
rect 5 -2356 7 -2344
rect 13 -2356 15 -2347
rect 56 -2356 58 -2334
rect -75 -2369 -73 -2366
rect -39 -2369 -37 -2366
rect -31 -2369 -29 -2366
rect 5 -2369 7 -2366
rect 13 -2369 15 -2366
rect 56 -2369 58 -2366
rect 835 -2367 837 -2364
rect 843 -2367 845 -2364
rect 873 -2367 875 -2364
rect 917 -2367 919 -2364
rect 962 -2367 964 -2364
rect 493 -2380 495 -2376
rect 195 -2417 197 -2414
rect 205 -2417 207 -2414
rect 606 -2381 608 -2377
rect 530 -2388 532 -2381
rect 563 -2395 565 -2381
rect 530 -2411 532 -2408
rect 563 -2418 565 -2415
rect 236 -2430 238 -2427
rect 195 -2462 197 -2441
rect 205 -2462 207 -2441
rect 493 -2440 495 -2420
rect 835 -2399 837 -2392
rect 830 -2403 837 -2399
rect 831 -2414 833 -2403
rect 843 -2411 845 -2392
rect 873 -2400 875 -2392
rect 917 -2400 919 -2392
rect 867 -2402 875 -2400
rect 911 -2402 919 -2400
rect 867 -2414 869 -2402
rect 875 -2414 877 -2405
rect 911 -2414 913 -2402
rect 919 -2414 921 -2405
rect 962 -2414 964 -2392
rect 530 -2428 532 -2425
rect 236 -2456 238 -2442
rect 563 -2435 565 -2432
rect 96 -2470 98 -2467
rect 106 -2470 108 -2467
rect 236 -2465 238 -2462
rect 493 -2463 495 -2460
rect 530 -2462 532 -2448
rect 606 -2441 608 -2421
rect 831 -2427 833 -2424
rect 867 -2427 869 -2424
rect 875 -2427 877 -2424
rect 911 -2427 913 -2424
rect 919 -2427 921 -2424
rect 962 -2427 964 -2424
rect 563 -2462 565 -2455
rect 606 -2464 608 -2461
rect 136 -2471 138 -2468
rect 195 -2471 197 -2468
rect 205 -2471 207 -2468
rect 96 -2502 98 -2482
rect 106 -2502 108 -2482
rect 136 -2497 138 -2483
rect 136 -2506 138 -2503
rect -834 -2518 -832 -2515
rect -826 -2518 -824 -2515
rect -796 -2518 -794 -2515
rect -752 -2518 -750 -2515
rect -707 -2518 -705 -2515
rect -621 -2518 -619 -2515
rect -613 -2518 -611 -2515
rect -583 -2518 -581 -2515
rect -539 -2518 -537 -2515
rect -494 -2518 -492 -2515
rect 96 -2517 98 -2514
rect 106 -2517 108 -2514
rect -128 -2538 -126 -2535
rect -118 -2538 -116 -2535
rect -834 -2550 -832 -2543
rect -839 -2554 -832 -2550
rect -838 -2565 -836 -2554
rect -826 -2562 -824 -2543
rect -796 -2551 -794 -2543
rect -752 -2551 -750 -2543
rect -802 -2553 -794 -2551
rect -758 -2553 -750 -2551
rect -802 -2565 -800 -2553
rect -794 -2565 -792 -2556
rect -758 -2565 -756 -2553
rect -750 -2565 -748 -2556
rect -707 -2565 -705 -2543
rect -621 -2550 -619 -2543
rect -626 -2554 -619 -2550
rect -625 -2565 -623 -2554
rect -613 -2562 -611 -2543
rect -583 -2551 -581 -2543
rect -539 -2551 -537 -2543
rect -589 -2553 -581 -2551
rect -545 -2553 -537 -2551
rect -589 -2565 -587 -2553
rect -581 -2565 -579 -2556
rect -545 -2565 -543 -2553
rect -537 -2565 -535 -2556
rect -494 -2565 -492 -2543
rect -374 -2549 -372 -2545
rect -838 -2578 -836 -2575
rect -802 -2578 -800 -2575
rect -794 -2578 -792 -2575
rect -758 -2578 -756 -2575
rect -750 -2578 -748 -2575
rect -707 -2578 -705 -2575
rect -625 -2578 -623 -2575
rect -589 -2578 -587 -2575
rect -581 -2578 -579 -2575
rect -545 -2578 -543 -2575
rect -537 -2578 -535 -2575
rect -494 -2578 -492 -2575
rect -261 -2550 -259 -2546
rect -88 -2539 -86 -2536
rect -337 -2557 -335 -2550
rect -304 -2564 -302 -2550
rect -337 -2580 -335 -2577
rect -304 -2587 -302 -2584
rect -374 -2609 -372 -2589
rect -128 -2570 -126 -2550
rect -118 -2570 -116 -2550
rect -88 -2565 -86 -2551
rect -88 -2574 -86 -2571
rect -128 -2585 -126 -2582
rect -118 -2585 -116 -2582
rect -337 -2597 -335 -2594
rect -304 -2604 -302 -2601
rect -374 -2632 -372 -2629
rect -337 -2631 -335 -2617
rect -261 -2610 -259 -2590
rect -304 -2631 -302 -2624
rect -261 -2633 -259 -2630
rect 825 -2675 827 -2672
rect 833 -2675 835 -2672
rect 863 -2675 865 -2672
rect 907 -2675 909 -2672
rect 952 -2675 954 -2672
rect 483 -2688 485 -2684
rect 103 -2713 105 -2710
rect 113 -2713 115 -2710
rect 143 -2714 145 -2711
rect 103 -2745 105 -2725
rect 113 -2745 115 -2725
rect 143 -2740 145 -2726
rect 596 -2689 598 -2685
rect 520 -2696 522 -2689
rect 553 -2703 555 -2689
rect 520 -2719 522 -2716
rect 553 -2726 555 -2723
rect 143 -2749 145 -2746
rect 483 -2748 485 -2728
rect 825 -2707 827 -2700
rect 820 -2711 827 -2707
rect 821 -2722 823 -2711
rect 833 -2719 835 -2700
rect 863 -2708 865 -2700
rect 907 -2708 909 -2700
rect 857 -2710 865 -2708
rect 901 -2710 909 -2708
rect 857 -2722 859 -2710
rect 865 -2722 867 -2713
rect 901 -2722 903 -2710
rect 909 -2722 911 -2713
rect 952 -2722 954 -2700
rect 520 -2736 522 -2733
rect 356 -2753 358 -2750
rect 366 -2753 368 -2750
rect 103 -2760 105 -2757
rect 113 -2760 115 -2757
rect 397 -2766 399 -2763
rect 205 -2782 207 -2779
rect 215 -2782 217 -2779
rect 246 -2795 248 -2792
rect 205 -2827 207 -2806
rect 215 -2827 217 -2806
rect 356 -2798 358 -2777
rect 366 -2798 368 -2777
rect 553 -2743 555 -2740
rect 483 -2771 485 -2768
rect 520 -2770 522 -2756
rect 596 -2749 598 -2729
rect 821 -2735 823 -2732
rect 857 -2735 859 -2732
rect 865 -2735 867 -2732
rect 901 -2735 903 -2732
rect 909 -2735 911 -2732
rect 952 -2735 954 -2732
rect 553 -2770 555 -2763
rect 596 -2772 598 -2769
rect 397 -2792 399 -2778
rect 397 -2801 399 -2798
rect 356 -2807 358 -2804
rect 366 -2807 368 -2804
rect 246 -2821 248 -2807
rect 106 -2835 108 -2832
rect 116 -2835 118 -2832
rect 246 -2830 248 -2827
rect -819 -2847 -817 -2844
rect -811 -2847 -809 -2844
rect -781 -2847 -779 -2844
rect -737 -2847 -735 -2844
rect -692 -2847 -690 -2844
rect -606 -2847 -604 -2844
rect -598 -2847 -596 -2844
rect -568 -2847 -566 -2844
rect -524 -2847 -522 -2844
rect -479 -2847 -477 -2844
rect 146 -2836 148 -2833
rect 205 -2836 207 -2833
rect 215 -2836 217 -2833
rect -113 -2867 -111 -2864
rect -103 -2867 -101 -2864
rect -819 -2879 -817 -2872
rect -824 -2883 -817 -2879
rect -823 -2894 -821 -2883
rect -811 -2891 -809 -2872
rect -781 -2880 -779 -2872
rect -737 -2880 -735 -2872
rect -787 -2882 -779 -2880
rect -743 -2882 -735 -2880
rect -787 -2894 -785 -2882
rect -779 -2894 -777 -2885
rect -743 -2894 -741 -2882
rect -735 -2894 -733 -2885
rect -692 -2894 -690 -2872
rect -606 -2879 -604 -2872
rect -611 -2883 -604 -2879
rect -610 -2894 -608 -2883
rect -598 -2891 -596 -2872
rect -568 -2880 -566 -2872
rect -524 -2880 -522 -2872
rect -574 -2882 -566 -2880
rect -530 -2882 -522 -2880
rect -574 -2894 -572 -2882
rect -566 -2894 -564 -2885
rect -530 -2894 -528 -2882
rect -522 -2894 -520 -2885
rect -479 -2894 -477 -2872
rect -359 -2878 -357 -2874
rect -823 -2907 -821 -2904
rect -787 -2907 -785 -2904
rect -779 -2907 -777 -2904
rect -743 -2907 -741 -2904
rect -735 -2907 -733 -2904
rect -692 -2907 -690 -2904
rect -610 -2907 -608 -2904
rect -574 -2907 -572 -2904
rect -566 -2907 -564 -2904
rect -530 -2907 -528 -2904
rect -522 -2907 -520 -2904
rect -479 -2907 -477 -2904
rect -246 -2879 -244 -2875
rect -73 -2868 -71 -2865
rect 106 -2867 108 -2847
rect 116 -2867 118 -2847
rect 146 -2862 148 -2848
rect -322 -2886 -320 -2879
rect -289 -2893 -287 -2879
rect -322 -2909 -320 -2906
rect -289 -2916 -287 -2913
rect -359 -2938 -357 -2918
rect -113 -2899 -111 -2879
rect -103 -2899 -101 -2879
rect 146 -2871 148 -2868
rect -73 -2894 -71 -2880
rect 106 -2882 108 -2879
rect 116 -2882 118 -2879
rect -73 -2903 -71 -2900
rect -113 -2914 -111 -2911
rect -103 -2914 -101 -2911
rect -322 -2926 -320 -2923
rect -289 -2933 -287 -2930
rect -359 -2961 -357 -2958
rect -322 -2960 -320 -2946
rect -246 -2939 -244 -2919
rect 849 -2934 851 -2931
rect 857 -2934 859 -2931
rect 887 -2934 889 -2931
rect 931 -2934 933 -2931
rect 976 -2934 978 -2931
rect -289 -2960 -287 -2953
rect 507 -2947 509 -2943
rect -246 -2962 -244 -2959
rect 101 -2977 103 -2974
rect 111 -2977 113 -2974
rect 141 -2978 143 -2975
rect 101 -3009 103 -2989
rect 111 -3009 113 -2989
rect 620 -2948 622 -2944
rect 544 -2955 546 -2948
rect 577 -2962 579 -2948
rect 544 -2978 546 -2975
rect 577 -2985 579 -2982
rect 141 -3004 143 -2990
rect 507 -3007 509 -2987
rect 849 -2966 851 -2959
rect 844 -2970 851 -2966
rect 845 -2981 847 -2970
rect 857 -2978 859 -2959
rect 887 -2967 889 -2959
rect 931 -2967 933 -2959
rect 881 -2969 889 -2967
rect 925 -2969 933 -2967
rect 881 -2981 883 -2969
rect 889 -2981 891 -2972
rect 925 -2981 927 -2969
rect 933 -2981 935 -2972
rect 976 -2981 978 -2959
rect 544 -2995 546 -2992
rect 141 -3013 143 -3010
rect 101 -3024 103 -3021
rect 111 -3024 113 -3021
rect 577 -3002 579 -2999
rect 507 -3030 509 -3027
rect 544 -3029 546 -3015
rect 620 -3008 622 -2988
rect 845 -2994 847 -2991
rect 881 -2994 883 -2991
rect 889 -2994 891 -2991
rect 925 -2994 927 -2991
rect 933 -2994 935 -2991
rect 976 -2994 978 -2991
rect 577 -3029 579 -3022
rect 620 -3031 622 -3028
rect 203 -3046 205 -3043
rect 213 -3046 215 -3043
rect 244 -3059 246 -3056
rect 203 -3091 205 -3070
rect 213 -3091 215 -3070
rect 244 -3085 246 -3071
rect 312 -3073 314 -3070
rect 322 -3073 324 -3070
rect 104 -3099 106 -3096
rect 114 -3099 116 -3096
rect 244 -3094 246 -3091
rect 353 -3086 355 -3083
rect 144 -3100 146 -3097
rect 203 -3100 205 -3097
rect 213 -3100 215 -3097
rect -795 -3114 -793 -3111
rect -787 -3114 -785 -3111
rect -757 -3114 -755 -3111
rect -713 -3114 -711 -3111
rect -668 -3114 -666 -3111
rect -582 -3114 -580 -3111
rect -574 -3114 -572 -3111
rect -544 -3114 -542 -3111
rect -500 -3114 -498 -3111
rect -455 -3114 -453 -3111
rect 104 -3131 106 -3111
rect 114 -3131 116 -3111
rect 144 -3126 146 -3112
rect 312 -3118 314 -3097
rect 322 -3118 324 -3097
rect 353 -3112 355 -3098
rect 353 -3121 355 -3118
rect -89 -3134 -87 -3131
rect -79 -3134 -77 -3131
rect -795 -3146 -793 -3139
rect -800 -3150 -793 -3146
rect -799 -3161 -797 -3150
rect -787 -3158 -785 -3139
rect -757 -3147 -755 -3139
rect -713 -3147 -711 -3139
rect -763 -3149 -755 -3147
rect -719 -3149 -711 -3147
rect -763 -3161 -761 -3149
rect -755 -3161 -753 -3152
rect -719 -3161 -717 -3149
rect -711 -3161 -709 -3152
rect -668 -3161 -666 -3139
rect -582 -3146 -580 -3139
rect -587 -3150 -580 -3146
rect -586 -3161 -584 -3150
rect -574 -3158 -572 -3139
rect -544 -3147 -542 -3139
rect -500 -3147 -498 -3139
rect -550 -3149 -542 -3147
rect -506 -3149 -498 -3147
rect -550 -3161 -548 -3149
rect -542 -3161 -540 -3152
rect -506 -3161 -504 -3149
rect -498 -3161 -496 -3152
rect -455 -3161 -453 -3139
rect -335 -3145 -333 -3141
rect -799 -3174 -797 -3171
rect -763 -3174 -761 -3171
rect -755 -3174 -753 -3171
rect -719 -3174 -717 -3171
rect -711 -3174 -709 -3171
rect -668 -3174 -666 -3171
rect -586 -3174 -584 -3171
rect -550 -3174 -548 -3171
rect -542 -3174 -540 -3171
rect -506 -3174 -504 -3171
rect -498 -3174 -496 -3171
rect -455 -3174 -453 -3171
rect -222 -3146 -220 -3142
rect -49 -3135 -47 -3132
rect -298 -3153 -296 -3146
rect -265 -3160 -263 -3146
rect -298 -3176 -296 -3173
rect -265 -3183 -263 -3180
rect -335 -3205 -333 -3185
rect -89 -3166 -87 -3146
rect -79 -3166 -77 -3146
rect 312 -3127 314 -3124
rect 322 -3127 324 -3124
rect 144 -3135 146 -3132
rect 205 -3133 207 -3130
rect 215 -3133 217 -3130
rect 104 -3146 106 -3143
rect 114 -3146 116 -3143
rect -49 -3161 -47 -3147
rect 246 -3146 248 -3143
rect -49 -3170 -47 -3167
rect 111 -3178 113 -3175
rect 121 -3178 123 -3175
rect -89 -3181 -87 -3178
rect -79 -3181 -77 -3178
rect -298 -3193 -296 -3190
rect -265 -3200 -263 -3197
rect -335 -3228 -333 -3225
rect -298 -3227 -296 -3213
rect -222 -3206 -220 -3186
rect 151 -3179 153 -3176
rect 205 -3178 207 -3157
rect 215 -3178 217 -3157
rect 246 -3172 248 -3158
rect -265 -3227 -263 -3220
rect 111 -3210 113 -3190
rect 121 -3210 123 -3190
rect 246 -3181 248 -3178
rect 205 -3187 207 -3184
rect 215 -3187 217 -3184
rect 151 -3205 153 -3191
rect 151 -3214 153 -3211
rect 111 -3225 113 -3222
rect 121 -3225 123 -3222
rect -222 -3229 -220 -3226
rect 870 -3240 872 -3237
rect 878 -3240 880 -3237
rect 908 -3240 910 -3237
rect 952 -3240 954 -3237
rect 997 -3240 999 -3237
rect 528 -3253 530 -3249
rect 641 -3254 643 -3250
rect 565 -3261 567 -3254
rect 598 -3268 600 -3254
rect 565 -3284 567 -3281
rect 598 -3291 600 -3288
rect 528 -3313 530 -3293
rect 870 -3272 872 -3265
rect 865 -3276 872 -3272
rect 866 -3287 868 -3276
rect 878 -3284 880 -3265
rect 908 -3273 910 -3265
rect 952 -3273 954 -3265
rect 902 -3275 910 -3273
rect 946 -3275 954 -3273
rect 902 -3287 904 -3275
rect 910 -3287 912 -3278
rect 946 -3287 948 -3275
rect 954 -3287 956 -3278
rect 997 -3287 999 -3265
rect 565 -3301 567 -3298
rect 107 -3322 109 -3319
rect 117 -3322 119 -3319
rect 147 -3323 149 -3320
rect 107 -3354 109 -3334
rect 117 -3354 119 -3334
rect 598 -3308 600 -3305
rect 147 -3349 149 -3335
rect 528 -3336 530 -3333
rect 565 -3335 567 -3321
rect 641 -3314 643 -3294
rect 866 -3300 868 -3297
rect 902 -3300 904 -3297
rect 910 -3300 912 -3297
rect 946 -3300 948 -3297
rect 954 -3300 956 -3297
rect 997 -3300 999 -3297
rect 598 -3335 600 -3328
rect 641 -3337 643 -3334
rect 147 -3358 149 -3355
rect 107 -3369 109 -3366
rect 117 -3369 119 -3366
rect 209 -3391 211 -3388
rect 219 -3391 221 -3388
rect 250 -3404 252 -3401
rect -766 -3424 -764 -3421
rect -758 -3424 -756 -3421
rect -728 -3424 -726 -3421
rect -684 -3424 -682 -3421
rect -639 -3424 -637 -3421
rect -553 -3424 -551 -3421
rect -545 -3424 -543 -3421
rect -515 -3424 -513 -3421
rect -471 -3424 -469 -3421
rect -426 -3424 -424 -3421
rect 209 -3436 211 -3415
rect 219 -3436 221 -3415
rect 250 -3430 252 -3416
rect 318 -3418 320 -3415
rect 328 -3418 330 -3415
rect -60 -3444 -58 -3441
rect -50 -3444 -48 -3441
rect -766 -3456 -764 -3449
rect -771 -3460 -764 -3456
rect -770 -3471 -768 -3460
rect -758 -3468 -756 -3449
rect -728 -3457 -726 -3449
rect -684 -3457 -682 -3449
rect -734 -3459 -726 -3457
rect -690 -3459 -682 -3457
rect -734 -3471 -732 -3459
rect -726 -3471 -724 -3462
rect -690 -3471 -688 -3459
rect -682 -3471 -680 -3462
rect -639 -3471 -637 -3449
rect -553 -3456 -551 -3449
rect -558 -3460 -551 -3456
rect -557 -3471 -555 -3460
rect -545 -3468 -543 -3449
rect -515 -3457 -513 -3449
rect -471 -3457 -469 -3449
rect -521 -3459 -513 -3457
rect -477 -3459 -469 -3457
rect -521 -3471 -519 -3459
rect -513 -3471 -511 -3462
rect -477 -3471 -475 -3459
rect -469 -3471 -467 -3462
rect -426 -3471 -424 -3449
rect -306 -3455 -304 -3451
rect -770 -3484 -768 -3481
rect -734 -3484 -732 -3481
rect -726 -3484 -724 -3481
rect -690 -3484 -688 -3481
rect -682 -3484 -680 -3481
rect -639 -3484 -637 -3481
rect -557 -3484 -555 -3481
rect -521 -3484 -519 -3481
rect -513 -3484 -511 -3481
rect -477 -3484 -475 -3481
rect -469 -3484 -467 -3481
rect -426 -3484 -424 -3481
rect -193 -3456 -191 -3452
rect -20 -3445 -18 -3442
rect 110 -3444 112 -3441
rect 120 -3444 122 -3441
rect 250 -3439 252 -3436
rect 359 -3431 361 -3428
rect -269 -3463 -267 -3456
rect -236 -3470 -234 -3456
rect -269 -3486 -267 -3483
rect -236 -3493 -234 -3490
rect -306 -3515 -304 -3495
rect -60 -3476 -58 -3456
rect -50 -3476 -48 -3456
rect 150 -3445 152 -3442
rect 209 -3445 211 -3442
rect 219 -3445 221 -3442
rect -20 -3471 -18 -3457
rect 110 -3476 112 -3456
rect 120 -3476 122 -3456
rect 150 -3471 152 -3457
rect 318 -3463 320 -3442
rect 328 -3463 330 -3442
rect 420 -3442 422 -3439
rect 430 -3442 432 -3439
rect 610 -3442 612 -3439
rect 618 -3442 620 -3439
rect 648 -3442 650 -3439
rect 692 -3442 694 -3439
rect 737 -3442 739 -3439
rect 359 -3457 361 -3443
rect 359 -3466 361 -3463
rect 461 -3455 463 -3452
rect -20 -3480 -18 -3477
rect 318 -3472 320 -3469
rect 328 -3472 330 -3469
rect 150 -3480 152 -3477
rect 211 -3478 213 -3475
rect 221 -3478 223 -3475
rect -60 -3491 -58 -3488
rect -50 -3491 -48 -3488
rect 110 -3491 112 -3488
rect 120 -3491 122 -3488
rect -269 -3503 -267 -3500
rect -236 -3510 -234 -3507
rect -306 -3538 -304 -3535
rect -269 -3537 -267 -3523
rect -193 -3516 -191 -3496
rect 420 -3487 422 -3466
rect 430 -3487 432 -3466
rect 461 -3481 463 -3467
rect 610 -3474 612 -3467
rect 605 -3478 612 -3474
rect 252 -3491 254 -3488
rect -236 -3537 -234 -3530
rect 117 -3523 119 -3520
rect 127 -3523 129 -3520
rect 157 -3524 159 -3521
rect 211 -3523 213 -3502
rect 221 -3523 223 -3502
rect 461 -3490 463 -3487
rect 606 -3489 608 -3478
rect 618 -3486 620 -3467
rect 648 -3475 650 -3467
rect 692 -3475 694 -3467
rect 642 -3477 650 -3475
rect 686 -3477 694 -3475
rect 642 -3489 644 -3477
rect 650 -3489 652 -3480
rect 686 -3489 688 -3477
rect 694 -3489 696 -3480
rect 737 -3489 739 -3467
rect 420 -3496 422 -3493
rect 430 -3496 432 -3493
rect 606 -3502 608 -3499
rect 642 -3502 644 -3499
rect 650 -3502 652 -3499
rect 686 -3502 688 -3499
rect 694 -3502 696 -3499
rect 737 -3502 739 -3499
rect 252 -3517 254 -3503
rect -193 -3539 -191 -3536
rect 117 -3555 119 -3535
rect 127 -3555 129 -3535
rect 252 -3526 254 -3523
rect 211 -3532 213 -3529
rect 221 -3532 223 -3529
rect 157 -3550 159 -3536
rect 157 -3559 159 -3556
rect 117 -3570 119 -3567
rect 127 -3570 129 -3567
rect 117 -3605 119 -3602
rect 127 -3605 129 -3602
rect 157 -3606 159 -3603
rect 117 -3637 119 -3617
rect 127 -3637 129 -3617
rect 157 -3632 159 -3618
rect 157 -3641 159 -3638
rect 117 -3652 119 -3649
rect 127 -3652 129 -3649
<< polycontact >>
rect -80 -2345 -76 -2341
rect -67 -2353 -63 -2349
rect -44 -2353 -39 -2348
rect -29 -2353 -24 -2349
rect 0 -2353 5 -2348
rect 52 -2348 56 -2343
rect 15 -2353 20 -2349
rect 529 -2381 533 -2376
rect 562 -2381 566 -2376
rect 191 -2459 195 -2455
rect 201 -2452 205 -2448
rect 489 -2437 493 -2432
rect 826 -2403 830 -2399
rect 839 -2411 843 -2407
rect 862 -2411 867 -2406
rect 877 -2411 882 -2407
rect 906 -2411 911 -2406
rect 958 -2406 962 -2401
rect 921 -2411 926 -2407
rect 232 -2453 236 -2449
rect 602 -2438 606 -2433
rect 529 -2467 533 -2462
rect 562 -2467 566 -2462
rect 92 -2493 96 -2489
rect 102 -2499 106 -2495
rect 132 -2494 136 -2490
rect -843 -2554 -839 -2550
rect -830 -2562 -826 -2558
rect -807 -2562 -802 -2557
rect -792 -2562 -787 -2558
rect -763 -2562 -758 -2557
rect -711 -2557 -707 -2552
rect -748 -2562 -743 -2558
rect -630 -2554 -626 -2550
rect -617 -2562 -613 -2558
rect -594 -2562 -589 -2557
rect -579 -2562 -574 -2558
rect -550 -2562 -545 -2557
rect -498 -2557 -494 -2552
rect -535 -2562 -530 -2558
rect -338 -2550 -334 -2545
rect -305 -2550 -301 -2545
rect -378 -2606 -374 -2601
rect -132 -2561 -128 -2557
rect -122 -2567 -118 -2563
rect -92 -2562 -88 -2558
rect -265 -2607 -261 -2602
rect -338 -2636 -334 -2631
rect -305 -2636 -301 -2631
rect 99 -2736 103 -2732
rect 109 -2742 113 -2738
rect 139 -2737 143 -2733
rect 519 -2689 523 -2684
rect 552 -2689 556 -2684
rect 479 -2745 483 -2740
rect 816 -2711 820 -2707
rect 829 -2719 833 -2715
rect 852 -2719 857 -2714
rect 867 -2719 872 -2715
rect 896 -2719 901 -2714
rect 948 -2714 952 -2709
rect 911 -2719 916 -2715
rect 352 -2795 356 -2791
rect 201 -2824 205 -2820
rect 211 -2817 215 -2813
rect 362 -2788 366 -2784
rect 592 -2746 596 -2741
rect 519 -2775 523 -2770
rect 552 -2775 556 -2770
rect 393 -2789 397 -2785
rect 242 -2818 246 -2814
rect 102 -2858 106 -2854
rect -828 -2883 -824 -2879
rect -815 -2891 -811 -2887
rect -792 -2891 -787 -2886
rect -777 -2891 -772 -2887
rect -748 -2891 -743 -2886
rect -696 -2886 -692 -2881
rect -733 -2891 -728 -2887
rect -615 -2883 -611 -2879
rect -602 -2891 -598 -2887
rect -579 -2891 -574 -2886
rect -564 -2891 -559 -2887
rect -535 -2891 -530 -2886
rect -483 -2886 -479 -2881
rect -520 -2891 -515 -2887
rect -323 -2879 -319 -2874
rect -290 -2879 -286 -2874
rect 112 -2864 116 -2860
rect 142 -2859 146 -2855
rect -363 -2935 -359 -2930
rect -117 -2890 -113 -2886
rect -107 -2896 -103 -2892
rect -77 -2891 -73 -2887
rect -250 -2936 -246 -2931
rect -323 -2965 -319 -2960
rect -290 -2965 -286 -2960
rect 97 -3000 101 -2996
rect 107 -3006 111 -3002
rect 543 -2948 547 -2943
rect 576 -2948 580 -2943
rect 137 -3001 141 -2997
rect 503 -3004 507 -2999
rect 840 -2970 844 -2966
rect 853 -2978 857 -2974
rect 876 -2978 881 -2973
rect 891 -2978 896 -2974
rect 920 -2978 925 -2973
rect 972 -2973 976 -2968
rect 935 -2978 940 -2974
rect 616 -3005 620 -3000
rect 543 -3034 547 -3029
rect 576 -3034 580 -3029
rect 199 -3088 203 -3084
rect 209 -3081 213 -3077
rect 240 -3082 244 -3078
rect 100 -3122 104 -3118
rect 110 -3128 114 -3124
rect 140 -3123 144 -3119
rect 308 -3115 312 -3111
rect 318 -3108 322 -3104
rect 349 -3109 353 -3105
rect -804 -3150 -800 -3146
rect -791 -3158 -787 -3154
rect -768 -3158 -763 -3153
rect -753 -3158 -748 -3154
rect -724 -3158 -719 -3153
rect -672 -3153 -668 -3148
rect -709 -3158 -704 -3154
rect -591 -3150 -587 -3146
rect -578 -3158 -574 -3154
rect -555 -3158 -550 -3153
rect -540 -3158 -535 -3154
rect -511 -3158 -506 -3153
rect -459 -3153 -455 -3148
rect -496 -3158 -491 -3154
rect -299 -3146 -295 -3141
rect -266 -3146 -262 -3141
rect -339 -3202 -335 -3197
rect -93 -3157 -89 -3153
rect -83 -3163 -79 -3159
rect -53 -3158 -49 -3154
rect 201 -3175 205 -3171
rect -226 -3203 -222 -3198
rect 211 -3168 215 -3164
rect 242 -3169 246 -3165
rect 107 -3201 111 -3197
rect 117 -3207 121 -3203
rect 147 -3202 151 -3198
rect -299 -3232 -295 -3227
rect -266 -3232 -262 -3227
rect 564 -3254 568 -3249
rect 597 -3254 601 -3249
rect 524 -3310 528 -3305
rect 861 -3276 865 -3272
rect 874 -3284 878 -3280
rect 897 -3284 902 -3279
rect 912 -3284 917 -3280
rect 941 -3284 946 -3279
rect 993 -3279 997 -3274
rect 956 -3284 961 -3280
rect 103 -3345 107 -3341
rect 113 -3351 117 -3347
rect 143 -3346 147 -3342
rect 637 -3311 641 -3306
rect 564 -3340 568 -3335
rect 597 -3340 601 -3335
rect 205 -3433 209 -3429
rect 215 -3426 219 -3422
rect 246 -3427 250 -3423
rect -775 -3460 -771 -3456
rect -762 -3468 -758 -3464
rect -739 -3468 -734 -3463
rect -724 -3468 -719 -3464
rect -695 -3468 -690 -3463
rect -643 -3463 -639 -3458
rect -680 -3468 -675 -3464
rect -562 -3460 -558 -3456
rect -549 -3468 -545 -3464
rect -526 -3468 -521 -3463
rect -511 -3468 -506 -3464
rect -482 -3468 -477 -3463
rect -430 -3463 -426 -3458
rect -467 -3468 -462 -3464
rect -270 -3456 -266 -3451
rect -237 -3456 -233 -3451
rect -310 -3512 -306 -3507
rect -64 -3467 -60 -3463
rect -54 -3473 -50 -3469
rect -24 -3468 -20 -3464
rect 106 -3467 110 -3463
rect 116 -3473 120 -3469
rect 146 -3468 150 -3464
rect 314 -3460 318 -3456
rect 324 -3453 328 -3449
rect 355 -3454 359 -3450
rect -197 -3513 -193 -3508
rect 416 -3484 420 -3480
rect 426 -3477 430 -3473
rect 457 -3478 461 -3474
rect 601 -3478 605 -3474
rect 207 -3520 211 -3516
rect 217 -3513 221 -3509
rect 614 -3486 618 -3482
rect 637 -3486 642 -3481
rect 652 -3486 657 -3482
rect 681 -3486 686 -3481
rect 733 -3481 737 -3476
rect 696 -3486 701 -3482
rect 248 -3514 252 -3510
rect -270 -3542 -266 -3537
rect -237 -3542 -233 -3537
rect 113 -3546 117 -3542
rect 123 -3552 127 -3548
rect 153 -3547 157 -3543
rect 113 -3628 117 -3624
rect 123 -3634 127 -3630
rect 153 -3629 157 -3625
<< metal1 >>
rect 317 -2299 324 -2298
rect -82 -2303 71 -2299
rect -76 -2309 -72 -2303
rect -38 -2309 -34 -2303
rect 6 -2309 10 -2303
rect 51 -2309 55 -2303
rect 317 -2308 705 -2299
rect -26 -2334 -13 -2309
rect 18 -2334 31 -2309
rect -87 -2345 -80 -2341
rect -60 -2342 -56 -2334
rect -60 -2345 -20 -2342
rect -70 -2353 -67 -2349
rect -60 -2356 -56 -2345
rect -48 -2353 -44 -2348
rect -24 -2353 -20 -2345
rect -16 -2348 -13 -2334
rect 28 -2343 31 -2334
rect 28 -2348 52 -2343
rect 59 -2344 63 -2334
rect 317 -2344 324 -2308
rect 460 -2344 685 -2339
rect 59 -2348 324 -2344
rect -16 -2353 0 -2348
rect 20 -2353 24 -2349
rect -16 -2356 -13 -2353
rect 28 -2356 31 -2348
rect 59 -2349 321 -2348
rect 59 -2356 63 -2349
rect -68 -2366 -56 -2356
rect -24 -2366 -13 -2356
rect 20 -2366 31 -2356
rect -80 -2371 -76 -2366
rect -44 -2371 -40 -2366
rect 0 -2371 4 -2366
rect 51 -2371 55 -2366
rect -81 -2375 63 -2371
rect 73 -2490 78 -2349
rect 488 -2380 492 -2344
rect 146 -2411 226 -2408
rect 85 -2462 128 -2461
rect 146 -2462 149 -2411
rect 190 -2417 193 -2411
rect 223 -2421 226 -2411
rect 513 -2412 518 -2357
rect 529 -2376 533 -2369
rect 562 -2376 566 -2369
rect 601 -2381 605 -2344
rect 698 -2358 705 -2308
rect 648 -2364 705 -2358
rect 824 -2361 977 -2357
rect 621 -2369 705 -2364
rect 830 -2367 834 -2361
rect 868 -2367 872 -2361
rect 912 -2367 916 -2361
rect 957 -2367 961 -2361
rect 525 -2412 529 -2408
rect 513 -2416 529 -2412
rect 223 -2424 249 -2421
rect 85 -2464 149 -2462
rect 91 -2470 94 -2464
rect 110 -2470 113 -2464
rect 125 -2465 149 -2464
rect 166 -2452 201 -2449
rect 209 -2450 212 -2441
rect 231 -2430 234 -2424
rect 479 -2437 489 -2432
rect 496 -2433 500 -2420
rect 525 -2428 529 -2416
rect 496 -2438 509 -2433
rect 496 -2440 500 -2438
rect 131 -2471 134 -2465
rect 100 -2485 103 -2482
rect 100 -2488 113 -2485
rect 73 -2493 92 -2490
rect 110 -2491 113 -2488
rect 110 -2494 132 -2491
rect 140 -2491 143 -2483
rect 166 -2491 171 -2452
rect 209 -2453 232 -2450
rect 240 -2450 243 -2442
rect 240 -2453 321 -2450
rect 174 -2458 191 -2455
rect 209 -2456 212 -2453
rect 240 -2456 243 -2453
rect 200 -2459 212 -2456
rect 200 -2462 203 -2459
rect 231 -2466 234 -2462
rect 190 -2474 193 -2468
rect 209 -2474 212 -2468
rect 221 -2469 249 -2466
rect 221 -2474 225 -2469
rect 140 -2494 171 -2491
rect 182 -2477 225 -2474
rect 45 -2499 102 -2496
rect 110 -2502 113 -2494
rect 140 -2497 143 -2494
rect -845 -2512 -141 -2508
rect -839 -2518 -835 -2512
rect -801 -2518 -797 -2512
rect -757 -2518 -753 -2512
rect -712 -2518 -708 -2512
rect -626 -2518 -622 -2512
rect -588 -2518 -584 -2512
rect -544 -2518 -540 -2512
rect -499 -2518 -495 -2512
rect -407 -2513 -141 -2512
rect -789 -2543 -776 -2518
rect -745 -2543 -732 -2518
rect -576 -2543 -563 -2518
rect -532 -2543 -519 -2518
rect -850 -2554 -843 -2550
rect -823 -2551 -819 -2543
rect -823 -2554 -783 -2551
rect -833 -2562 -830 -2558
rect -823 -2565 -819 -2554
rect -811 -2562 -807 -2557
rect -787 -2562 -783 -2554
rect -779 -2557 -776 -2543
rect -735 -2552 -732 -2543
rect -735 -2557 -711 -2552
rect -704 -2553 -700 -2543
rect -779 -2562 -763 -2557
rect -743 -2562 -739 -2558
rect -779 -2565 -776 -2562
rect -735 -2565 -732 -2557
rect -704 -2558 -691 -2553
rect -704 -2565 -700 -2558
rect -637 -2554 -630 -2550
rect -610 -2551 -606 -2543
rect -610 -2554 -570 -2551
rect -620 -2562 -617 -2558
rect -610 -2565 -606 -2554
rect -598 -2562 -594 -2557
rect -574 -2562 -570 -2554
rect -566 -2557 -563 -2543
rect -522 -2552 -519 -2543
rect -522 -2557 -498 -2552
rect -491 -2553 -487 -2543
rect -379 -2549 -375 -2513
rect -566 -2562 -550 -2557
rect -530 -2562 -526 -2558
rect -566 -2565 -563 -2562
rect -522 -2565 -519 -2557
rect -491 -2558 -478 -2553
rect -491 -2565 -487 -2558
rect -831 -2575 -819 -2565
rect -787 -2575 -776 -2565
rect -743 -2575 -732 -2565
rect -618 -2575 -606 -2565
rect -574 -2575 -563 -2565
rect -530 -2575 -519 -2565
rect -843 -2580 -839 -2575
rect -807 -2580 -803 -2575
rect -763 -2580 -759 -2575
rect -712 -2580 -708 -2575
rect -630 -2580 -626 -2575
rect -594 -2580 -590 -2575
rect -550 -2580 -546 -2575
rect -499 -2580 -495 -2575
rect -844 -2584 -487 -2580
rect -491 -2669 -487 -2584
rect -354 -2581 -349 -2526
rect -338 -2545 -334 -2538
rect -305 -2545 -301 -2538
rect -266 -2550 -262 -2513
rect -179 -2533 -173 -2526
rect -146 -2529 -141 -2513
rect 131 -2507 134 -2503
rect 182 -2507 186 -2477
rect 121 -2510 186 -2507
rect 91 -2520 94 -2514
rect 121 -2520 125 -2510
rect 85 -2523 125 -2520
rect -146 -2530 -96 -2529
rect -146 -2532 -75 -2530
rect -246 -2538 -165 -2533
rect -342 -2581 -338 -2577
rect -354 -2585 -338 -2581
rect -388 -2606 -378 -2601
rect -371 -2602 -367 -2589
rect -342 -2597 -338 -2585
rect -371 -2607 -358 -2602
rect -371 -2609 -367 -2607
rect -334 -2582 -330 -2577
rect -334 -2586 -317 -2582
rect -334 -2597 -330 -2586
rect -321 -2596 -317 -2586
rect -309 -2596 -305 -2584
rect -321 -2601 -305 -2596
rect -379 -2668 -375 -2629
rect -338 -2649 -334 -2636
rect -321 -2660 -315 -2601
rect -309 -2604 -305 -2601
rect -301 -2597 -297 -2584
rect -301 -2601 -280 -2597
rect -301 -2604 -297 -2601
rect -286 -2602 -280 -2601
rect -286 -2607 -276 -2602
rect -270 -2607 -265 -2602
rect -258 -2603 -254 -2590
rect -216 -2564 -207 -2551
rect -168 -2558 -165 -2538
rect -133 -2538 -130 -2532
rect -114 -2538 -111 -2532
rect -99 -2533 -75 -2532
rect -93 -2539 -90 -2533
rect -124 -2553 -121 -2550
rect -124 -2556 -111 -2553
rect -168 -2561 -132 -2558
rect -114 -2559 -111 -2556
rect -114 -2562 -92 -2559
rect -84 -2559 -81 -2551
rect -84 -2562 -33 -2559
rect -216 -2567 -122 -2564
rect -258 -2608 -241 -2603
rect -258 -2610 -254 -2608
rect -305 -2649 -301 -2636
rect -266 -2668 -262 -2630
rect -216 -2648 -208 -2567
rect -114 -2570 -111 -2562
rect -84 -2565 -81 -2562
rect -93 -2575 -90 -2571
rect -103 -2578 -75 -2575
rect -133 -2588 -130 -2582
rect -103 -2588 -99 -2578
rect -198 -2591 -99 -2588
rect -198 -2668 -187 -2591
rect 317 -2630 321 -2453
rect 533 -2413 537 -2408
rect 533 -2417 550 -2413
rect 533 -2428 537 -2417
rect 546 -2427 550 -2417
rect 558 -2427 562 -2415
rect 546 -2432 562 -2427
rect 488 -2499 492 -2460
rect 529 -2480 533 -2467
rect 546 -2490 552 -2432
rect 558 -2435 562 -2432
rect 566 -2428 570 -2415
rect 880 -2392 893 -2367
rect 924 -2392 937 -2367
rect 809 -2403 826 -2399
rect 846 -2400 850 -2392
rect 846 -2403 886 -2400
rect 836 -2411 839 -2407
rect 846 -2414 850 -2403
rect 858 -2411 862 -2406
rect 882 -2411 886 -2403
rect 890 -2406 893 -2392
rect 934 -2401 937 -2392
rect 934 -2406 958 -2401
rect 965 -2402 969 -2392
rect 890 -2411 906 -2406
rect 926 -2411 930 -2407
rect 890 -2414 893 -2411
rect 934 -2414 937 -2406
rect 965 -2407 978 -2402
rect 965 -2414 969 -2407
rect 566 -2432 587 -2428
rect 566 -2435 570 -2432
rect 581 -2433 587 -2432
rect 581 -2438 591 -2433
rect 597 -2438 602 -2433
rect 609 -2434 613 -2421
rect 838 -2424 850 -2414
rect 882 -2424 893 -2414
rect 926 -2424 937 -2414
rect 826 -2429 830 -2424
rect 862 -2429 866 -2424
rect 906 -2429 910 -2424
rect 957 -2429 961 -2424
rect 825 -2433 969 -2429
rect 609 -2439 626 -2434
rect 609 -2441 613 -2439
rect 651 -2442 722 -2436
rect 562 -2480 566 -2467
rect 601 -2499 605 -2461
rect 651 -2479 659 -2442
rect 460 -2507 669 -2499
rect 706 -2589 722 -2442
rect 705 -2630 715 -2629
rect 317 -2636 715 -2630
rect 450 -2652 683 -2647
rect -407 -2669 -187 -2668
rect -491 -2676 -187 -2669
rect 478 -2688 482 -2652
rect 92 -2705 135 -2704
rect 155 -2705 198 -2704
rect 92 -2707 198 -2705
rect 98 -2713 101 -2707
rect 117 -2713 120 -2707
rect 132 -2708 198 -2707
rect 138 -2714 141 -2708
rect 107 -2728 110 -2725
rect 107 -2731 120 -2728
rect -18 -2736 99 -2733
rect 117 -2734 120 -2731
rect -830 -2841 -126 -2837
rect -824 -2847 -820 -2841
rect -786 -2847 -782 -2841
rect -742 -2847 -738 -2841
rect -697 -2847 -693 -2841
rect -611 -2847 -607 -2841
rect -573 -2847 -569 -2841
rect -529 -2847 -525 -2841
rect -484 -2847 -480 -2841
rect -392 -2842 -126 -2841
rect -774 -2872 -761 -2847
rect -730 -2872 -717 -2847
rect -561 -2872 -548 -2847
rect -517 -2872 -504 -2847
rect -835 -2883 -828 -2879
rect -808 -2880 -804 -2872
rect -808 -2883 -768 -2880
rect -818 -2891 -815 -2887
rect -808 -2894 -804 -2883
rect -796 -2891 -792 -2886
rect -772 -2891 -768 -2883
rect -764 -2886 -761 -2872
rect -720 -2881 -717 -2872
rect -720 -2886 -696 -2881
rect -689 -2882 -685 -2872
rect -764 -2891 -748 -2886
rect -728 -2891 -724 -2887
rect -764 -2894 -761 -2891
rect -720 -2894 -717 -2886
rect -689 -2887 -676 -2882
rect -689 -2894 -685 -2887
rect -622 -2883 -615 -2879
rect -595 -2880 -591 -2872
rect -595 -2883 -555 -2880
rect -605 -2891 -602 -2887
rect -595 -2894 -591 -2883
rect -583 -2891 -579 -2886
rect -559 -2891 -555 -2883
rect -551 -2886 -548 -2872
rect -507 -2881 -504 -2872
rect -507 -2886 -483 -2881
rect -476 -2882 -472 -2872
rect -364 -2878 -360 -2842
rect -551 -2891 -535 -2886
rect -515 -2891 -511 -2887
rect -551 -2894 -548 -2891
rect -507 -2894 -504 -2886
rect -476 -2887 -463 -2882
rect -476 -2894 -472 -2887
rect -816 -2904 -804 -2894
rect -772 -2904 -761 -2894
rect -728 -2904 -717 -2894
rect -603 -2904 -591 -2894
rect -559 -2904 -548 -2894
rect -515 -2904 -504 -2894
rect -828 -2909 -824 -2904
rect -792 -2909 -788 -2904
rect -748 -2909 -744 -2904
rect -697 -2909 -693 -2904
rect -615 -2909 -611 -2904
rect -579 -2909 -575 -2904
rect -535 -2909 -531 -2904
rect -484 -2909 -480 -2904
rect -829 -2913 -472 -2909
rect -476 -2998 -472 -2913
rect -339 -2910 -334 -2855
rect -323 -2874 -319 -2867
rect -290 -2874 -286 -2867
rect -251 -2879 -247 -2842
rect -164 -2862 -158 -2855
rect -131 -2858 -126 -2842
rect -18 -2855 -11 -2736
rect 117 -2737 139 -2734
rect 147 -2734 150 -2726
rect 147 -2737 167 -2734
rect 66 -2742 109 -2739
rect 117 -2745 120 -2737
rect 147 -2740 150 -2737
rect 138 -2750 141 -2746
rect 128 -2753 156 -2750
rect 98 -2763 101 -2757
rect 128 -2763 132 -2753
rect 92 -2766 132 -2763
rect 194 -2773 198 -2708
rect 503 -2720 508 -2665
rect 519 -2684 523 -2677
rect 552 -2684 556 -2677
rect 591 -2689 595 -2652
rect 638 -2667 689 -2666
rect 705 -2667 715 -2636
rect 638 -2672 715 -2667
rect 814 -2669 967 -2665
rect 611 -2677 715 -2672
rect 683 -2678 715 -2677
rect 820 -2675 824 -2669
rect 858 -2675 862 -2669
rect 902 -2675 906 -2669
rect 947 -2675 951 -2669
rect 515 -2720 519 -2716
rect 503 -2724 519 -2720
rect 257 -2744 346 -2743
rect 257 -2747 387 -2744
rect 469 -2745 479 -2740
rect 486 -2741 490 -2728
rect 515 -2736 519 -2724
rect 194 -2776 236 -2773
rect 200 -2782 203 -2776
rect 233 -2786 236 -2776
rect 257 -2785 260 -2747
rect 351 -2753 354 -2747
rect 384 -2757 387 -2747
rect 486 -2746 499 -2741
rect 486 -2748 490 -2746
rect 384 -2760 410 -2757
rect 256 -2786 260 -2785
rect 233 -2788 260 -2786
rect 295 -2788 362 -2785
rect 370 -2786 373 -2777
rect 392 -2766 395 -2760
rect 233 -2789 259 -2788
rect 175 -2817 211 -2814
rect 219 -2815 222 -2806
rect 241 -2795 244 -2789
rect 95 -2827 138 -2826
rect 95 -2829 159 -2827
rect 101 -2835 104 -2829
rect 120 -2835 123 -2829
rect 135 -2830 159 -2829
rect 141 -2836 144 -2830
rect 110 -2850 113 -2847
rect 110 -2853 123 -2850
rect -18 -2858 102 -2855
rect 120 -2856 123 -2853
rect -131 -2859 -81 -2858
rect -131 -2861 -60 -2859
rect -231 -2867 -150 -2862
rect -327 -2910 -323 -2906
rect -339 -2914 -323 -2910
rect -373 -2935 -363 -2930
rect -356 -2931 -352 -2918
rect -327 -2926 -323 -2914
rect -356 -2936 -343 -2931
rect -356 -2938 -352 -2936
rect -319 -2911 -315 -2906
rect -319 -2915 -302 -2911
rect -319 -2926 -315 -2915
rect -306 -2925 -302 -2915
rect -294 -2925 -290 -2913
rect -306 -2930 -290 -2925
rect -364 -2997 -360 -2958
rect -323 -2978 -319 -2965
rect -306 -2987 -300 -2930
rect -294 -2933 -290 -2930
rect -286 -2926 -282 -2913
rect -286 -2930 -265 -2926
rect -286 -2933 -282 -2930
rect -271 -2931 -265 -2930
rect -271 -2936 -261 -2931
rect -255 -2936 -250 -2931
rect -243 -2932 -239 -2919
rect -201 -2893 -192 -2880
rect -153 -2887 -150 -2867
rect -118 -2867 -115 -2861
rect -99 -2867 -96 -2861
rect -84 -2862 -60 -2861
rect -78 -2868 -75 -2862
rect -109 -2882 -106 -2879
rect -109 -2885 -96 -2882
rect -153 -2890 -117 -2887
rect -99 -2888 -96 -2885
rect -99 -2891 -77 -2888
rect -69 -2888 -66 -2880
rect -69 -2891 -46 -2888
rect -201 -2896 -107 -2893
rect -243 -2937 -226 -2932
rect -243 -2939 -239 -2937
rect -290 -2978 -286 -2965
rect -251 -2997 -247 -2959
rect -201 -2977 -193 -2896
rect -99 -2899 -96 -2891
rect -69 -2894 -66 -2891
rect -57 -2892 -46 -2891
rect -78 -2904 -75 -2900
rect -88 -2907 -60 -2904
rect -118 -2917 -115 -2911
rect -88 -2917 -84 -2907
rect -183 -2920 -84 -2917
rect -183 -2997 -172 -2920
rect -18 -2931 -11 -2858
rect 120 -2859 142 -2856
rect 150 -2856 153 -2848
rect 175 -2856 178 -2817
rect 219 -2818 242 -2815
rect 250 -2815 253 -2807
rect 295 -2815 299 -2788
rect 370 -2789 393 -2786
rect 401 -2786 404 -2778
rect 523 -2721 527 -2716
rect 523 -2725 540 -2721
rect 523 -2736 527 -2725
rect 536 -2735 540 -2725
rect 548 -2735 552 -2723
rect 536 -2740 552 -2735
rect 401 -2789 424 -2786
rect 330 -2794 352 -2791
rect 370 -2792 373 -2789
rect 401 -2792 404 -2789
rect 361 -2795 373 -2792
rect 361 -2798 364 -2795
rect 392 -2802 395 -2798
rect 351 -2810 354 -2804
rect 370 -2810 373 -2804
rect 382 -2805 410 -2802
rect 382 -2810 386 -2805
rect 250 -2818 299 -2815
rect 339 -2813 386 -2810
rect 184 -2823 201 -2820
rect 184 -2832 188 -2823
rect 219 -2821 222 -2818
rect 250 -2821 253 -2818
rect 210 -2824 222 -2821
rect 210 -2827 213 -2824
rect 241 -2831 244 -2827
rect 339 -2831 342 -2813
rect 200 -2839 203 -2833
rect 219 -2839 222 -2833
rect 231 -2834 322 -2831
rect 325 -2834 342 -2831
rect 231 -2839 235 -2834
rect 150 -2859 178 -2856
rect 190 -2842 235 -2839
rect -5 -2864 112 -2861
rect -5 -2865 7 -2864
rect 120 -2867 123 -2859
rect 150 -2862 153 -2859
rect 141 -2872 144 -2868
rect 190 -2872 194 -2842
rect 131 -2875 194 -2872
rect 101 -2885 104 -2879
rect 131 -2885 135 -2875
rect 95 -2888 135 -2885
rect 264 -2931 268 -2858
rect 419 -2879 424 -2789
rect 478 -2807 482 -2768
rect 519 -2788 523 -2775
rect 536 -2798 542 -2740
rect 548 -2743 552 -2740
rect 556 -2736 560 -2723
rect 870 -2700 883 -2675
rect 914 -2700 927 -2675
rect 799 -2711 816 -2707
rect 836 -2708 840 -2700
rect 836 -2711 876 -2708
rect 826 -2719 829 -2715
rect 836 -2722 840 -2711
rect 848 -2719 852 -2714
rect 872 -2719 876 -2711
rect 880 -2714 883 -2700
rect 924 -2709 927 -2700
rect 924 -2714 948 -2709
rect 955 -2710 959 -2700
rect 880 -2719 896 -2714
rect 916 -2719 920 -2715
rect 880 -2722 883 -2719
rect 924 -2722 927 -2714
rect 955 -2715 968 -2710
rect 955 -2722 959 -2715
rect 556 -2740 577 -2736
rect 556 -2743 560 -2740
rect 571 -2741 577 -2740
rect 571 -2746 581 -2741
rect 587 -2746 592 -2741
rect 599 -2742 603 -2729
rect 828 -2732 840 -2722
rect 872 -2732 883 -2722
rect 916 -2732 927 -2722
rect 816 -2737 820 -2732
rect 852 -2737 856 -2732
rect 896 -2737 900 -2732
rect 947 -2737 951 -2732
rect 815 -2741 959 -2737
rect 599 -2747 616 -2742
rect 599 -2749 603 -2747
rect 641 -2750 741 -2744
rect 552 -2788 556 -2775
rect 591 -2807 595 -2769
rect 641 -2787 649 -2750
rect 450 -2815 659 -2807
rect 419 -2885 722 -2879
rect 474 -2911 707 -2906
rect -19 -2935 268 -2931
rect -18 -2987 -11 -2935
rect 502 -2947 506 -2911
rect 90 -2969 133 -2968
rect 90 -2971 154 -2969
rect -105 -2993 -11 -2987
rect 96 -2977 99 -2971
rect 115 -2977 118 -2971
rect 130 -2972 154 -2971
rect 136 -2978 139 -2972
rect -392 -2998 -172 -2997
rect -476 -3005 -172 -2998
rect 105 -2992 108 -2989
rect 527 -2979 532 -2924
rect 543 -2943 547 -2936
rect 576 -2943 580 -2936
rect 615 -2948 619 -2911
rect 712 -2925 722 -2885
rect 662 -2931 722 -2925
rect 838 -2928 991 -2924
rect 635 -2936 722 -2931
rect 844 -2934 848 -2928
rect 882 -2934 886 -2928
rect 926 -2934 930 -2928
rect 971 -2934 975 -2928
rect 539 -2979 543 -2975
rect 527 -2983 543 -2979
rect 105 -2995 118 -2992
rect 52 -3000 97 -2997
rect 115 -2998 118 -2995
rect 115 -3001 137 -2998
rect 145 -2998 148 -2990
rect 145 -3001 165 -2998
rect 72 -3006 107 -3003
rect 115 -3009 118 -3001
rect 145 -3004 148 -3001
rect 136 -3014 139 -3010
rect 126 -3017 154 -3014
rect 96 -3027 99 -3021
rect 126 -3027 130 -3017
rect 90 -3030 130 -3027
rect 162 -3078 165 -3001
rect 493 -3004 503 -2999
rect 510 -3000 514 -2987
rect 539 -2995 543 -2983
rect 510 -3005 523 -3000
rect 510 -3007 514 -3005
rect 547 -2980 551 -2975
rect 547 -2984 564 -2980
rect 547 -2995 551 -2984
rect 560 -2994 564 -2984
rect 572 -2994 576 -2982
rect 560 -2999 576 -2994
rect 192 -3040 234 -3037
rect 198 -3046 201 -3040
rect 231 -3050 234 -3040
rect 231 -3053 257 -3050
rect 162 -3081 209 -3078
rect 217 -3079 220 -3070
rect 239 -3059 242 -3053
rect 301 -3067 343 -3064
rect 502 -3066 506 -3027
rect 543 -3047 547 -3034
rect 560 -3057 566 -2999
rect 572 -3002 576 -2999
rect 580 -2995 584 -2982
rect 894 -2959 907 -2934
rect 938 -2959 951 -2934
rect 823 -2970 840 -2966
rect 860 -2967 864 -2959
rect 860 -2970 900 -2967
rect 850 -2978 853 -2974
rect 860 -2981 864 -2970
rect 872 -2978 876 -2973
rect 896 -2978 900 -2970
rect 904 -2973 907 -2959
rect 948 -2968 951 -2959
rect 948 -2973 972 -2968
rect 979 -2969 983 -2959
rect 904 -2978 920 -2973
rect 940 -2978 944 -2974
rect 904 -2981 907 -2978
rect 948 -2981 951 -2973
rect 979 -2974 992 -2969
rect 979 -2981 983 -2974
rect 580 -2999 601 -2995
rect 580 -3002 584 -2999
rect 595 -3000 601 -2999
rect 595 -3005 605 -3000
rect 611 -3005 616 -3000
rect 623 -3001 627 -2988
rect 852 -2991 864 -2981
rect 896 -2991 907 -2981
rect 940 -2991 951 -2981
rect 840 -2996 844 -2991
rect 876 -2996 880 -2991
rect 920 -2996 924 -2991
rect 971 -2996 975 -2991
rect 839 -3000 983 -2996
rect 623 -3006 640 -3001
rect 704 -3003 713 -3002
rect 623 -3008 627 -3006
rect 665 -3009 715 -3003
rect 576 -3047 580 -3034
rect 615 -3066 619 -3028
rect 665 -3046 673 -3009
rect 217 -3082 240 -3079
rect 248 -3079 251 -3071
rect 307 -3073 310 -3067
rect 248 -3082 270 -3079
rect 173 -3087 199 -3084
rect 217 -3085 220 -3082
rect 248 -3085 251 -3082
rect 208 -3088 220 -3085
rect 93 -3091 136 -3090
rect 208 -3091 211 -3088
rect 93 -3093 157 -3091
rect 99 -3099 102 -3093
rect 118 -3099 121 -3093
rect 133 -3094 157 -3093
rect -806 -3108 -102 -3104
rect -800 -3114 -796 -3108
rect -762 -3114 -758 -3108
rect -718 -3114 -714 -3108
rect -673 -3114 -669 -3108
rect -587 -3114 -583 -3108
rect -549 -3114 -545 -3108
rect -505 -3114 -501 -3108
rect -460 -3114 -456 -3108
rect -368 -3109 -102 -3108
rect -750 -3139 -737 -3114
rect -706 -3139 -693 -3114
rect -537 -3139 -524 -3114
rect -493 -3139 -480 -3114
rect -811 -3150 -804 -3146
rect -784 -3147 -780 -3139
rect -784 -3150 -744 -3147
rect -794 -3158 -791 -3154
rect -784 -3161 -780 -3150
rect -772 -3158 -768 -3153
rect -748 -3158 -744 -3150
rect -740 -3153 -737 -3139
rect -696 -3148 -693 -3139
rect -696 -3153 -672 -3148
rect -665 -3149 -661 -3139
rect -740 -3158 -724 -3153
rect -704 -3158 -700 -3154
rect -740 -3161 -737 -3158
rect -696 -3161 -693 -3153
rect -665 -3154 -652 -3149
rect -665 -3161 -661 -3154
rect -598 -3150 -591 -3146
rect -571 -3147 -567 -3139
rect -571 -3150 -531 -3147
rect -581 -3158 -578 -3154
rect -571 -3161 -567 -3150
rect -559 -3158 -555 -3153
rect -535 -3158 -531 -3150
rect -527 -3153 -524 -3139
rect -483 -3148 -480 -3139
rect -483 -3153 -459 -3148
rect -452 -3149 -448 -3139
rect -340 -3145 -336 -3109
rect -527 -3158 -511 -3153
rect -491 -3158 -487 -3154
rect -527 -3161 -524 -3158
rect -483 -3161 -480 -3153
rect -452 -3154 -439 -3149
rect -452 -3161 -448 -3154
rect -792 -3171 -780 -3161
rect -748 -3171 -737 -3161
rect -704 -3171 -693 -3161
rect -579 -3171 -567 -3161
rect -535 -3171 -524 -3161
rect -491 -3171 -480 -3161
rect -804 -3176 -800 -3171
rect -768 -3176 -764 -3171
rect -724 -3176 -720 -3171
rect -673 -3176 -669 -3171
rect -591 -3176 -587 -3171
rect -555 -3176 -551 -3171
rect -511 -3176 -507 -3171
rect -460 -3176 -456 -3171
rect -805 -3180 -448 -3176
rect -452 -3265 -448 -3180
rect -315 -3177 -310 -3122
rect -299 -3141 -295 -3134
rect -266 -3141 -262 -3134
rect -227 -3146 -223 -3109
rect -140 -3129 -134 -3122
rect -107 -3125 -102 -3109
rect 139 -3100 142 -3094
rect 239 -3095 242 -3091
rect 108 -3114 111 -3111
rect 198 -3103 201 -3097
rect 217 -3103 220 -3097
rect 229 -3098 257 -3095
rect 229 -3103 233 -3098
rect 192 -3106 233 -3103
rect 267 -3105 270 -3082
rect 340 -3077 343 -3067
rect 474 -3074 683 -3066
rect 704 -3073 714 -3009
rect 340 -3080 366 -3077
rect 267 -3108 318 -3105
rect 326 -3106 329 -3097
rect 348 -3086 351 -3080
rect 326 -3109 349 -3106
rect 357 -3106 360 -3098
rect 705 -3100 714 -3099
rect 357 -3109 744 -3106
rect 108 -3117 121 -3114
rect 17 -3119 23 -3117
rect 17 -3122 100 -3119
rect 118 -3120 121 -3117
rect 118 -3123 140 -3120
rect 148 -3120 151 -3112
rect 264 -3114 308 -3111
rect 148 -3123 168 -3120
rect -107 -3126 -57 -3125
rect -107 -3128 -36 -3126
rect -207 -3134 -126 -3129
rect -303 -3177 -299 -3173
rect -315 -3181 -299 -3177
rect -349 -3202 -339 -3197
rect -332 -3198 -328 -3185
rect -303 -3193 -299 -3181
rect -332 -3203 -319 -3198
rect -332 -3205 -328 -3203
rect -295 -3178 -291 -3173
rect -295 -3182 -278 -3178
rect -295 -3193 -291 -3182
rect -282 -3192 -278 -3182
rect -270 -3192 -266 -3180
rect -282 -3197 -266 -3192
rect -340 -3264 -336 -3225
rect -299 -3245 -295 -3232
rect -282 -3258 -276 -3197
rect -270 -3200 -266 -3197
rect -262 -3193 -258 -3180
rect -262 -3197 -241 -3193
rect -262 -3200 -258 -3197
rect -247 -3198 -241 -3197
rect -247 -3203 -237 -3198
rect -231 -3203 -226 -3198
rect -219 -3199 -215 -3186
rect -177 -3160 -168 -3147
rect -129 -3154 -126 -3134
rect -94 -3134 -91 -3128
rect -75 -3134 -72 -3128
rect -60 -3129 -36 -3128
rect 86 -3128 110 -3125
rect -54 -3135 -51 -3129
rect -85 -3149 -82 -3146
rect -85 -3152 -72 -3149
rect -129 -3157 -93 -3154
rect -75 -3155 -72 -3152
rect -75 -3158 -53 -3155
rect -45 -3155 -42 -3147
rect -45 -3158 -24 -3155
rect -177 -3163 -83 -3160
rect -219 -3204 -202 -3199
rect -219 -3206 -215 -3204
rect -266 -3245 -262 -3232
rect -227 -3264 -223 -3226
rect -177 -3244 -169 -3163
rect -75 -3166 -72 -3158
rect -45 -3161 -42 -3158
rect -54 -3171 -51 -3167
rect -64 -3174 -36 -3171
rect -94 -3184 -91 -3178
rect -64 -3184 -60 -3174
rect -159 -3187 -60 -3184
rect -159 -3264 -148 -3187
rect 86 -3198 90 -3128
rect 118 -3131 121 -3123
rect 148 -3126 151 -3123
rect 139 -3136 142 -3132
rect 129 -3139 157 -3136
rect 99 -3149 102 -3143
rect 129 -3149 133 -3139
rect 93 -3152 133 -3149
rect 165 -3164 168 -3123
rect 194 -3127 236 -3124
rect 200 -3133 203 -3127
rect 233 -3137 236 -3127
rect 233 -3140 259 -3137
rect 165 -3165 170 -3164
rect 165 -3167 211 -3165
rect 167 -3168 211 -3167
rect 219 -3166 222 -3157
rect 241 -3146 244 -3140
rect 219 -3169 242 -3166
rect 250 -3166 253 -3158
rect 264 -3166 267 -3114
rect 326 -3112 329 -3109
rect 357 -3112 360 -3109
rect 317 -3115 329 -3112
rect 317 -3118 320 -3115
rect 348 -3122 351 -3118
rect 307 -3130 310 -3124
rect 326 -3130 329 -3124
rect 338 -3125 366 -3122
rect 338 -3130 342 -3125
rect 301 -3133 342 -3130
rect 250 -3169 267 -3166
rect 371 -3165 695 -3153
rect 100 -3170 143 -3169
rect 100 -3172 164 -3170
rect 106 -3178 109 -3172
rect 125 -3178 128 -3172
rect 140 -3173 164 -3172
rect 146 -3179 149 -3173
rect 181 -3174 201 -3171
rect 115 -3193 118 -3190
rect 115 -3196 128 -3193
rect 86 -3201 107 -3198
rect 125 -3199 128 -3196
rect 125 -3202 147 -3199
rect 155 -3199 158 -3191
rect 181 -3199 185 -3174
rect 219 -3172 222 -3169
rect 250 -3172 253 -3169
rect 210 -3175 222 -3172
rect 210 -3178 213 -3175
rect 241 -3182 244 -3178
rect 200 -3190 203 -3184
rect 219 -3190 222 -3184
rect 231 -3185 259 -3182
rect 231 -3190 235 -3185
rect 194 -3193 235 -3190
rect 155 -3202 185 -3199
rect -6 -3207 117 -3204
rect 125 -3210 128 -3202
rect 155 -3205 158 -3202
rect 146 -3215 149 -3211
rect 136 -3218 164 -3215
rect 106 -3228 109 -3222
rect 136 -3228 140 -3218
rect 100 -3231 140 -3228
rect -368 -3265 -148 -3264
rect -452 -3272 -148 -3265
rect -76 -3282 -60 -3253
rect 371 -3282 382 -3165
rect 738 -3212 744 -3109
rect 495 -3217 728 -3212
rect -77 -3295 382 -3282
rect 523 -3253 527 -3217
rect 548 -3285 553 -3230
rect 564 -3249 568 -3242
rect 597 -3249 601 -3242
rect 636 -3254 640 -3217
rect 738 -3231 743 -3212
rect 683 -3237 743 -3231
rect 859 -3234 1012 -3230
rect 656 -3241 743 -3237
rect 865 -3240 869 -3234
rect 903 -3240 907 -3234
rect 947 -3240 951 -3234
rect 992 -3240 996 -3234
rect 656 -3242 742 -3241
rect 729 -3243 742 -3242
rect 560 -3285 564 -3281
rect 548 -3289 564 -3285
rect -75 -3296 382 -3295
rect 514 -3310 524 -3305
rect 531 -3306 535 -3293
rect 560 -3301 564 -3289
rect 531 -3311 544 -3306
rect 531 -3313 535 -3311
rect 96 -3314 139 -3313
rect 96 -3316 160 -3314
rect 102 -3322 105 -3316
rect 121 -3322 124 -3316
rect 136 -3317 160 -3316
rect 142 -3323 145 -3317
rect 111 -3337 114 -3334
rect 111 -3340 124 -3337
rect 44 -3345 103 -3342
rect 121 -3343 124 -3340
rect 121 -3346 143 -3343
rect 151 -3343 154 -3335
rect 568 -3286 572 -3281
rect 568 -3290 585 -3286
rect 568 -3301 572 -3290
rect 581 -3300 585 -3290
rect 593 -3300 597 -3288
rect 581 -3305 597 -3300
rect 151 -3346 404 -3343
rect 93 -3351 113 -3348
rect 121 -3354 124 -3346
rect 151 -3349 154 -3346
rect 230 -3347 404 -3346
rect 396 -3353 404 -3347
rect 142 -3359 145 -3355
rect 132 -3362 160 -3359
rect 102 -3372 105 -3366
rect 132 -3372 136 -3362
rect 523 -3372 527 -3333
rect 564 -3353 568 -3340
rect 581 -3363 587 -3305
rect 593 -3308 597 -3305
rect 601 -3301 605 -3288
rect 915 -3265 928 -3240
rect 959 -3265 972 -3240
rect 844 -3276 861 -3272
rect 881 -3273 885 -3265
rect 881 -3276 921 -3273
rect 871 -3284 874 -3280
rect 881 -3287 885 -3276
rect 893 -3284 897 -3279
rect 917 -3284 921 -3276
rect 925 -3279 928 -3265
rect 969 -3274 972 -3265
rect 969 -3279 993 -3274
rect 1000 -3275 1004 -3265
rect 925 -3284 941 -3279
rect 961 -3284 965 -3280
rect 925 -3287 928 -3284
rect 969 -3287 972 -3279
rect 1000 -3280 1013 -3275
rect 1000 -3287 1004 -3280
rect 601 -3305 622 -3301
rect 601 -3308 605 -3305
rect 616 -3306 622 -3305
rect 616 -3311 626 -3306
rect 632 -3311 637 -3306
rect 644 -3307 648 -3294
rect 873 -3297 885 -3287
rect 917 -3297 928 -3287
rect 961 -3297 972 -3287
rect 861 -3302 865 -3297
rect 897 -3302 901 -3297
rect 941 -3302 945 -3297
rect 992 -3302 996 -3297
rect 860 -3306 1004 -3302
rect 644 -3312 661 -3307
rect 644 -3314 648 -3312
rect 686 -3315 725 -3309
rect 597 -3353 601 -3340
rect 636 -3372 640 -3334
rect 686 -3352 694 -3315
rect 96 -3375 136 -3372
rect 495 -3380 704 -3372
rect 198 -3385 240 -3382
rect 204 -3391 207 -3385
rect -231 -3414 -73 -3413
rect -777 -3418 -73 -3414
rect 237 -3395 240 -3385
rect 237 -3398 263 -3395
rect -771 -3424 -767 -3418
rect -733 -3424 -729 -3418
rect -689 -3424 -685 -3418
rect -644 -3424 -640 -3418
rect -558 -3424 -554 -3418
rect -520 -3424 -516 -3418
rect -476 -3424 -472 -3418
rect -431 -3424 -427 -3418
rect -339 -3419 -73 -3418
rect -721 -3449 -708 -3424
rect -677 -3449 -664 -3424
rect -508 -3449 -495 -3424
rect -464 -3449 -451 -3424
rect -782 -3460 -775 -3456
rect -755 -3457 -751 -3449
rect -755 -3460 -715 -3457
rect -765 -3468 -762 -3464
rect -755 -3471 -751 -3460
rect -743 -3468 -739 -3463
rect -719 -3468 -715 -3460
rect -711 -3463 -708 -3449
rect -667 -3458 -664 -3449
rect -667 -3463 -643 -3458
rect -636 -3459 -632 -3449
rect -711 -3468 -695 -3463
rect -675 -3468 -671 -3464
rect -711 -3471 -708 -3468
rect -667 -3471 -664 -3463
rect -636 -3464 -623 -3459
rect -636 -3471 -632 -3464
rect -569 -3460 -562 -3456
rect -542 -3457 -538 -3449
rect -542 -3460 -502 -3457
rect -552 -3468 -549 -3464
rect -542 -3471 -538 -3460
rect -530 -3468 -526 -3463
rect -506 -3468 -502 -3460
rect -498 -3463 -495 -3449
rect -454 -3458 -451 -3449
rect -454 -3463 -430 -3458
rect -423 -3459 -419 -3449
rect -311 -3455 -307 -3419
rect -231 -3420 -73 -3419
rect -498 -3468 -482 -3463
rect -462 -3468 -458 -3464
rect -498 -3471 -495 -3468
rect -454 -3471 -451 -3463
rect -423 -3464 -410 -3459
rect -423 -3471 -419 -3464
rect -763 -3481 -751 -3471
rect -719 -3481 -708 -3471
rect -675 -3481 -664 -3471
rect -550 -3481 -538 -3471
rect -506 -3481 -495 -3471
rect -462 -3481 -451 -3471
rect -775 -3486 -771 -3481
rect -739 -3486 -735 -3481
rect -695 -3486 -691 -3481
rect -644 -3486 -640 -3481
rect -562 -3486 -558 -3481
rect -526 -3486 -522 -3481
rect -482 -3486 -478 -3481
rect -431 -3486 -427 -3481
rect -776 -3490 -419 -3486
rect -423 -3575 -419 -3490
rect -286 -3487 -281 -3432
rect -270 -3451 -266 -3444
rect -237 -3451 -233 -3444
rect -198 -3456 -194 -3420
rect -111 -3439 -105 -3432
rect -78 -3435 -73 -3420
rect 38 -3426 215 -3423
rect 223 -3424 226 -3415
rect 245 -3404 248 -3398
rect 713 -3402 724 -3315
rect 307 -3412 349 -3409
rect -78 -3436 -28 -3435
rect -78 -3438 -7 -3436
rect -178 -3444 -97 -3439
rect -274 -3487 -270 -3483
rect -286 -3491 -270 -3487
rect -320 -3512 -310 -3507
rect -303 -3508 -299 -3495
rect -274 -3503 -270 -3491
rect -303 -3513 -290 -3508
rect -303 -3515 -299 -3513
rect -266 -3488 -262 -3483
rect -266 -3492 -249 -3488
rect -266 -3503 -262 -3492
rect -253 -3502 -249 -3492
rect -241 -3502 -237 -3490
rect -253 -3507 -237 -3502
rect -311 -3574 -307 -3535
rect -270 -3555 -266 -3542
rect -253 -3564 -247 -3507
rect -241 -3510 -237 -3507
rect -233 -3503 -229 -3490
rect -233 -3507 -212 -3503
rect -233 -3510 -229 -3507
rect -218 -3508 -212 -3507
rect -218 -3513 -208 -3508
rect -202 -3513 -197 -3508
rect -190 -3509 -186 -3496
rect -148 -3470 -139 -3457
rect -100 -3464 -97 -3444
rect -65 -3444 -62 -3438
rect -46 -3444 -43 -3438
rect -31 -3439 -7 -3438
rect -25 -3445 -22 -3439
rect -56 -3459 -53 -3456
rect -56 -3462 -43 -3459
rect -100 -3467 -64 -3464
rect -46 -3465 -43 -3462
rect -46 -3468 -24 -3465
rect -16 -3465 -13 -3457
rect 38 -3465 44 -3426
rect 223 -3427 246 -3424
rect 254 -3424 257 -3416
rect 313 -3418 316 -3412
rect 254 -3427 275 -3424
rect 186 -3432 205 -3429
rect 99 -3436 142 -3435
rect 99 -3438 163 -3436
rect 105 -3444 108 -3438
rect 124 -3444 127 -3438
rect 139 -3439 163 -3438
rect 145 -3445 148 -3439
rect 114 -3459 117 -3456
rect -16 -3468 44 -3465
rect 114 -3462 127 -3459
rect 56 -3467 106 -3464
rect 124 -3465 127 -3462
rect 124 -3468 146 -3465
rect 154 -3465 157 -3457
rect 186 -3465 189 -3432
rect 223 -3430 226 -3427
rect 254 -3430 257 -3427
rect 214 -3433 226 -3430
rect 214 -3436 217 -3433
rect 245 -3440 248 -3436
rect 204 -3448 207 -3442
rect 223 -3448 226 -3442
rect 235 -3443 263 -3440
rect 235 -3448 239 -3443
rect 198 -3451 239 -3448
rect 271 -3450 275 -3427
rect 346 -3422 349 -3412
rect 346 -3425 372 -3422
rect 271 -3453 324 -3450
rect 332 -3451 335 -3442
rect 354 -3431 357 -3425
rect 409 -3436 451 -3433
rect 599 -3436 752 -3432
rect 332 -3454 355 -3451
rect 363 -3451 366 -3443
rect 415 -3442 418 -3436
rect 363 -3454 381 -3451
rect 154 -3468 189 -3465
rect 294 -3459 314 -3456
rect -148 -3473 -54 -3470
rect -190 -3514 -173 -3509
rect -190 -3516 -186 -3514
rect -237 -3555 -233 -3542
rect -198 -3574 -194 -3536
rect -148 -3554 -140 -3473
rect -46 -3476 -43 -3468
rect -16 -3471 -13 -3468
rect -5 -3469 43 -3468
rect 94 -3473 116 -3470
rect 124 -3476 127 -3468
rect 154 -3471 157 -3468
rect -25 -3481 -22 -3477
rect -35 -3484 -7 -3481
rect -65 -3494 -62 -3488
rect -35 -3494 -31 -3484
rect 200 -3472 242 -3469
rect 145 -3481 148 -3477
rect 206 -3478 209 -3472
rect 135 -3484 163 -3481
rect 105 -3494 108 -3488
rect 135 -3494 139 -3484
rect -130 -3497 -31 -3494
rect 99 -3497 139 -3494
rect -130 -3574 -119 -3497
rect 239 -3482 242 -3472
rect 239 -3485 265 -3482
rect 174 -3513 217 -3510
rect 225 -3511 228 -3502
rect 247 -3491 250 -3485
rect 106 -3515 149 -3514
rect 106 -3517 170 -3515
rect 112 -3523 115 -3517
rect 131 -3523 134 -3517
rect 146 -3518 170 -3517
rect 152 -3524 155 -3518
rect 121 -3538 124 -3535
rect 121 -3541 134 -3538
rect 97 -3546 113 -3543
rect 131 -3544 134 -3541
rect 131 -3547 153 -3544
rect 161 -3544 164 -3536
rect 174 -3544 177 -3513
rect 225 -3514 248 -3511
rect 256 -3511 259 -3503
rect 294 -3511 298 -3459
rect 332 -3457 335 -3454
rect 363 -3457 366 -3454
rect 323 -3460 335 -3457
rect 323 -3463 326 -3460
rect 354 -3467 357 -3463
rect 313 -3475 316 -3469
rect 332 -3475 335 -3469
rect 344 -3470 372 -3467
rect 344 -3475 348 -3470
rect 307 -3478 348 -3475
rect 378 -3474 381 -3454
rect 448 -3446 451 -3436
rect 605 -3442 609 -3436
rect 643 -3442 647 -3436
rect 687 -3442 691 -3436
rect 732 -3442 736 -3436
rect 448 -3449 474 -3446
rect 378 -3477 426 -3474
rect 434 -3475 437 -3466
rect 456 -3455 459 -3449
rect 655 -3467 668 -3442
rect 699 -3467 712 -3442
rect 434 -3478 457 -3475
rect 465 -3475 468 -3467
rect 587 -3475 601 -3474
rect 465 -3478 601 -3475
rect 621 -3475 625 -3467
rect 621 -3478 661 -3475
rect 401 -3483 416 -3480
rect 434 -3481 437 -3478
rect 465 -3481 468 -3478
rect 425 -3484 437 -3481
rect 425 -3487 428 -3484
rect 611 -3486 614 -3482
rect 456 -3491 459 -3487
rect 621 -3489 625 -3478
rect 633 -3486 637 -3481
rect 657 -3486 661 -3478
rect 665 -3481 668 -3467
rect 709 -3476 712 -3467
rect 709 -3481 733 -3476
rect 740 -3477 744 -3467
rect 665 -3486 681 -3481
rect 701 -3486 705 -3482
rect 665 -3489 668 -3486
rect 709 -3489 712 -3481
rect 740 -3482 753 -3477
rect 740 -3489 744 -3482
rect 415 -3499 418 -3493
rect 434 -3499 437 -3493
rect 446 -3494 474 -3491
rect 446 -3499 450 -3494
rect 409 -3502 450 -3499
rect 613 -3499 625 -3489
rect 657 -3499 668 -3489
rect 701 -3499 712 -3489
rect 601 -3504 605 -3499
rect 637 -3504 641 -3499
rect 681 -3504 685 -3499
rect 732 -3504 736 -3499
rect 600 -3508 744 -3504
rect 256 -3514 298 -3511
rect 161 -3547 177 -3544
rect 181 -3519 207 -3516
rect 84 -3552 123 -3549
rect 131 -3555 134 -3547
rect 161 -3550 164 -3547
rect 152 -3560 155 -3556
rect 142 -3563 170 -3560
rect 112 -3573 115 -3567
rect 142 -3573 146 -3563
rect -339 -3575 -119 -3574
rect -423 -3582 -119 -3575
rect 106 -3576 146 -3573
rect 106 -3597 149 -3596
rect 106 -3599 170 -3597
rect 112 -3605 115 -3599
rect 131 -3605 134 -3599
rect 146 -3600 170 -3599
rect 152 -3606 155 -3600
rect 121 -3620 124 -3617
rect 121 -3623 134 -3620
rect 91 -3628 113 -3625
rect 131 -3626 134 -3623
rect 131 -3629 153 -3626
rect 161 -3626 164 -3618
rect 181 -3626 185 -3519
rect 225 -3517 228 -3514
rect 256 -3517 259 -3514
rect 216 -3520 228 -3517
rect 216 -3523 219 -3520
rect 247 -3527 250 -3523
rect 206 -3535 209 -3529
rect 225 -3535 228 -3529
rect 237 -3530 265 -3527
rect 237 -3535 241 -3530
rect 200 -3538 241 -3535
rect 161 -3627 185 -3626
rect 161 -3629 184 -3627
rect 0 -3634 123 -3631
rect 131 -3637 134 -3629
rect 161 -3632 164 -3629
rect 152 -3642 155 -3638
rect 142 -3645 170 -3642
rect 112 -3655 115 -3649
rect 142 -3655 146 -3645
rect 106 -3658 146 -3655
<< m2contact >>
rect 513 -2357 519 -2352
rect 529 -2369 534 -2364
rect 561 -2369 566 -2364
rect 613 -2369 621 -2364
rect 474 -2437 479 -2432
rect 509 -2438 515 -2433
rect -691 -2559 -680 -2552
rect -354 -2526 -348 -2521
rect -478 -2559 -467 -2552
rect -338 -2538 -333 -2533
rect -306 -2538 -301 -2533
rect -182 -2526 -172 -2519
rect 151 -2499 158 -2494
rect -254 -2538 -246 -2533
rect -393 -2606 -388 -2601
rect -358 -2607 -352 -2602
rect -338 -2654 -333 -2649
rect -217 -2551 -206 -2545
rect -276 -2607 -270 -2602
rect -241 -2608 -235 -2603
rect -305 -2654 -300 -2649
rect -216 -2654 -208 -2648
rect 529 -2485 534 -2480
rect 804 -2404 809 -2399
rect 591 -2438 597 -2433
rect 626 -2439 632 -2434
rect 562 -2485 567 -2480
rect 546 -2496 552 -2490
rect 651 -2485 659 -2479
rect 503 -2665 509 -2660
rect -676 -2888 -665 -2881
rect -339 -2855 -333 -2850
rect -463 -2888 -452 -2881
rect -323 -2867 -318 -2862
rect -291 -2867 -286 -2862
rect -167 -2855 -157 -2848
rect 58 -2745 66 -2739
rect 163 -2742 168 -2737
rect 519 -2677 524 -2672
rect 551 -2677 556 -2672
rect 603 -2677 611 -2672
rect 464 -2745 469 -2740
rect 499 -2746 505 -2741
rect -239 -2867 -231 -2862
rect -378 -2935 -373 -2930
rect -343 -2936 -337 -2931
rect -323 -2983 -318 -2978
rect -202 -2880 -191 -2874
rect -261 -2936 -255 -2931
rect -226 -2937 -220 -2932
rect -290 -2983 -285 -2978
rect -306 -2992 -300 -2987
rect -201 -2983 -193 -2977
rect 325 -2796 330 -2791
rect 519 -2793 524 -2788
rect 794 -2712 799 -2707
rect 581 -2746 587 -2741
rect 616 -2747 622 -2742
rect 552 -2793 557 -2788
rect 536 -2804 542 -2798
rect 641 -2793 649 -2787
rect -113 -2993 -105 -2984
rect 527 -2924 533 -2919
rect 41 -3000 52 -2991
rect 543 -2936 548 -2931
rect 575 -2936 580 -2931
rect 627 -2936 635 -2931
rect 488 -3004 493 -2999
rect 523 -3005 529 -3000
rect 543 -3052 548 -3047
rect 818 -2971 823 -2966
rect 605 -3005 611 -3000
rect 640 -3006 646 -3001
rect 576 -3052 581 -3047
rect 560 -3063 566 -3057
rect 665 -3052 673 -3046
rect 162 -3086 167 -3081
rect -652 -3155 -641 -3148
rect -315 -3122 -309 -3117
rect -439 -3155 -428 -3148
rect -299 -3134 -294 -3129
rect -267 -3134 -262 -3129
rect -143 -3122 -133 -3115
rect 696 -3099 720 -3073
rect -215 -3134 -207 -3129
rect -354 -3202 -349 -3197
rect -319 -3203 -313 -3198
rect -299 -3250 -294 -3245
rect -178 -3147 -167 -3141
rect -237 -3203 -231 -3198
rect -202 -3204 -196 -3199
rect -266 -3250 -261 -3245
rect -177 -3250 -169 -3244
rect 158 -3167 165 -3161
rect 695 -3171 719 -3145
rect 548 -3230 554 -3225
rect 564 -3242 569 -3237
rect 596 -3242 601 -3237
rect 648 -3242 656 -3237
rect 509 -3310 514 -3305
rect 544 -3311 550 -3306
rect 32 -3346 44 -3337
rect 87 -3353 93 -3348
rect 396 -3362 404 -3353
rect 564 -3358 569 -3353
rect 839 -3277 844 -3272
rect 626 -3311 632 -3306
rect 661 -3312 667 -3307
rect 597 -3358 602 -3353
rect 581 -3369 587 -3363
rect 686 -3358 694 -3352
rect -623 -3465 -612 -3458
rect -286 -3432 -280 -3427
rect -410 -3465 -399 -3458
rect -270 -3444 -265 -3439
rect -238 -3444 -233 -3439
rect -114 -3432 -104 -3425
rect -186 -3444 -178 -3439
rect -325 -3512 -320 -3507
rect -290 -3513 -284 -3508
rect -270 -3560 -265 -3555
rect -149 -3457 -138 -3451
rect -208 -3513 -202 -3508
rect 56 -3464 62 -3459
rect 708 -3420 724 -3402
rect -173 -3514 -167 -3509
rect -237 -3560 -232 -3555
rect -254 -3570 -244 -3564
rect 87 -3475 94 -3470
rect -148 -3560 -140 -3554
rect 88 -3546 97 -3539
rect 396 -3485 401 -3480
rect 81 -3628 91 -3619
<< metal2 >>
rect 519 -2357 632 -2352
rect 474 -2369 529 -2364
rect 534 -2369 561 -2364
rect 566 -2369 613 -2364
rect 474 -2432 478 -2369
rect 509 -2480 515 -2438
rect 591 -2479 597 -2438
rect 626 -2434 632 -2357
rect 508 -2485 529 -2480
rect 534 -2485 562 -2480
rect 567 -2485 581 -2480
rect 591 -2485 651 -2479
rect -452 -2490 -448 -2489
rect -452 -2494 -174 -2490
rect -665 -2505 -470 -2501
rect -665 -2553 -661 -2505
rect -680 -2558 -661 -2553
rect -452 -2553 -448 -2494
rect -409 -2503 -209 -2499
rect -348 -2526 -235 -2521
rect -467 -2558 -448 -2553
rect -393 -2538 -338 -2533
rect -333 -2538 -306 -2533
rect -301 -2538 -254 -2533
rect -393 -2601 -389 -2538
rect -358 -2649 -352 -2607
rect -276 -2648 -270 -2607
rect -241 -2603 -235 -2526
rect -215 -2545 -209 -2503
rect -179 -2505 -174 -2494
rect 804 -2492 809 -2404
rect 552 -2496 809 -2492
rect -179 -2515 -173 -2505
rect -179 -2519 -174 -2515
rect -359 -2654 -338 -2649
rect -333 -2654 -305 -2649
rect -300 -2654 -286 -2649
rect -276 -2654 -216 -2648
rect 151 -2671 155 -2499
rect 509 -2665 622 -2660
rect 58 -2675 155 -2671
rect 58 -2739 62 -2675
rect 464 -2677 519 -2672
rect 524 -2677 551 -2672
rect 556 -2677 603 -2672
rect 464 -2740 468 -2677
rect 163 -2791 167 -2742
rect 499 -2788 505 -2746
rect 581 -2787 587 -2746
rect 616 -2742 622 -2665
rect 34 -2795 167 -2791
rect -437 -2819 -433 -2818
rect -437 -2823 -159 -2819
rect -650 -2834 -455 -2830
rect -650 -2882 -646 -2834
rect -665 -2887 -646 -2882
rect -437 -2882 -433 -2823
rect -394 -2832 -194 -2828
rect -333 -2855 -220 -2850
rect -452 -2887 -433 -2882
rect -378 -2867 -323 -2862
rect -318 -2867 -291 -2862
rect -286 -2867 -239 -2862
rect -378 -2930 -374 -2867
rect -343 -2978 -337 -2936
rect -261 -2977 -255 -2936
rect -226 -2932 -220 -2855
rect -200 -2874 -194 -2832
rect -164 -2834 -159 -2823
rect -164 -2848 -158 -2834
rect -344 -2983 -323 -2978
rect -318 -2983 -290 -2978
rect -285 -2983 -271 -2978
rect -261 -2983 -201 -2977
rect -300 -2992 -113 -2988
rect 34 -3000 41 -2795
rect 163 -2893 167 -2795
rect 322 -2893 325 -2791
rect 498 -2793 519 -2788
rect 524 -2793 552 -2788
rect 557 -2793 571 -2788
rect 581 -2793 641 -2787
rect 794 -2800 799 -2712
rect 542 -2804 799 -2800
rect 163 -2898 326 -2893
rect 533 -2924 646 -2919
rect 488 -2936 543 -2931
rect 548 -2936 575 -2931
rect 580 -2936 627 -2931
rect 488 -2999 492 -2936
rect 523 -3047 529 -3005
rect 605 -3046 611 -3005
rect 640 -3001 646 -2924
rect 522 -3052 543 -3047
rect 548 -3052 576 -3047
rect 581 -3052 595 -3047
rect 605 -3052 665 -3046
rect 818 -3059 823 -2971
rect 566 -3063 823 -3059
rect -413 -3086 -409 -3085
rect 32 -3086 162 -3081
rect -413 -3090 -135 -3086
rect -626 -3101 -431 -3097
rect -626 -3149 -622 -3101
rect -641 -3154 -622 -3149
rect -413 -3149 -409 -3090
rect -370 -3099 -170 -3095
rect -176 -3103 -170 -3099
rect -177 -3113 -170 -3103
rect -309 -3122 -196 -3117
rect -428 -3154 -409 -3149
rect -354 -3134 -299 -3129
rect -294 -3134 -267 -3129
rect -262 -3134 -215 -3129
rect -354 -3197 -350 -3134
rect -319 -3245 -313 -3203
rect -237 -3244 -231 -3203
rect -202 -3199 -196 -3122
rect -176 -3141 -170 -3113
rect -140 -3102 -135 -3090
rect -140 -3115 -134 -3102
rect -320 -3250 -299 -3245
rect -294 -3250 -266 -3245
rect -261 -3250 -247 -3245
rect -237 -3250 -177 -3244
rect 32 -3337 39 -3086
rect 703 -3115 716 -3099
rect 703 -3145 715 -3115
rect 56 -3165 158 -3161
rect -384 -3396 -380 -3395
rect -384 -3400 -106 -3396
rect -597 -3411 -402 -3407
rect -597 -3459 -593 -3411
rect -612 -3464 -593 -3459
rect -384 -3459 -380 -3400
rect -341 -3409 -141 -3405
rect -280 -3432 -167 -3427
rect -399 -3464 -380 -3459
rect -325 -3444 -270 -3439
rect -265 -3444 -238 -3439
rect -233 -3444 -186 -3439
rect -325 -3507 -321 -3444
rect -290 -3555 -284 -3513
rect -208 -3554 -202 -3513
rect -173 -3509 -167 -3432
rect -147 -3451 -141 -3409
rect -111 -3425 -106 -3400
rect 56 -3459 62 -3165
rect 554 -3230 667 -3225
rect 509 -3242 564 -3237
rect 569 -3242 596 -3237
rect 601 -3242 648 -3237
rect 509 -3305 513 -3242
rect 544 -3353 550 -3311
rect 626 -3352 632 -3311
rect 661 -3307 667 -3230
rect 88 -3470 93 -3353
rect 543 -3358 564 -3353
rect 569 -3358 597 -3353
rect 602 -3358 616 -3353
rect 626 -3358 686 -3352
rect 89 -3539 92 -3475
rect 396 -3480 401 -3362
rect 839 -3365 844 -3277
rect 587 -3369 844 -3365
rect 688 -3410 708 -3409
rect 544 -3412 708 -3410
rect 543 -3420 708 -3412
rect -291 -3560 -270 -3555
rect -265 -3560 -237 -3555
rect -232 -3560 -218 -3555
rect -208 -3560 -148 -3554
rect 89 -3566 92 -3546
rect -244 -3570 92 -3566
rect 83 -3583 88 -3570
rect 543 -3583 556 -3420
rect 83 -3592 556 -3583
rect 83 -3619 88 -3592
<< m3contact >>
rect -470 -2506 -457 -2500
rect -419 -2505 -409 -2499
rect 45 -2503 53 -2496
rect -321 -2665 -315 -2659
rect 706 -2589 730 -2572
rect 722 -2760 741 -2740
rect -455 -2835 -442 -2829
rect -404 -2834 -394 -2828
rect 172 -2864 178 -2859
rect 264 -2867 277 -2858
rect 72 -3008 78 -3003
rect -431 -3102 -418 -3096
rect -380 -3101 -370 -3095
rect 14 -3117 23 -3109
rect -282 -3259 -275 -3254
rect -75 -3270 -60 -3253
rect 82 -3130 90 -3125
rect -402 -3412 -389 -3406
rect -351 -3411 -341 -3405
rect 86 -3202 91 -3197
rect 167 -3207 172 -3202
rect 76 -3553 84 -3548
<< metal3 >>
rect -457 -2505 -419 -2500
rect 45 -2655 51 -2503
rect 327 -2581 706 -2578
rect 326 -2589 706 -2581
rect 326 -2590 726 -2589
rect 326 -2655 338 -2590
rect -321 -2659 338 -2655
rect -315 -2665 338 -2659
rect -442 -2834 -404 -2829
rect 173 -2949 178 -2864
rect 727 -2860 740 -2760
rect 277 -2867 740 -2860
rect 727 -2868 740 -2867
rect 14 -2958 178 -2949
rect -418 -3101 -380 -3096
rect 14 -3109 23 -2958
rect 72 -3125 76 -3008
rect 72 -3129 82 -3125
rect -275 -3258 -75 -3254
rect -60 -3255 44 -3254
rect 86 -3255 89 -3202
rect -60 -3258 92 -3255
rect 168 -3275 172 -3207
rect 76 -3279 172 -3275
rect -389 -3411 -351 -3406
rect 76 -3548 80 -3279
<< m4contact >>
rect 174 -2461 181 -2455
rect -36 -2565 -27 -2556
rect 183 -2832 190 -2827
rect -5 -2872 7 -2861
rect -57 -2896 -45 -2886
rect 173 -3089 181 -3084
rect -33 -3160 -24 -3153
rect -7 -3213 12 -3199
rect 0 -3639 10 -3629
<< metal4 >>
rect 159 -2442 165 -2441
rect -36 -2446 165 -2442
rect -36 -2556 -30 -2446
rect 159 -2455 165 -2446
rect 159 -2461 174 -2455
rect -27 -2565 5 -2561
rect -35 -2566 5 -2565
rect -5 -2861 3 -2566
rect -56 -2909 -49 -2896
rect -5 -2909 3 -2907
rect 184 -2909 187 -2832
rect -56 -2915 187 -2909
rect -32 -3250 -25 -3160
rect -5 -3199 3 -2915
rect 0 -3250 6 -3249
rect 174 -3250 178 -3089
rect -32 -3256 178 -3250
rect 0 -3629 6 -3256
<< labels >>
rlabel metal1 -77 -2562 -72 -2559 1 g0
rlabel metal1 -620 -2561 -618 -2559 1 clk
rlabel metal1 -597 -2561 -596 -2559 1 clk
rlabel metal1 -529 -2561 -527 -2559 1 clk
rlabel metal1 -485 -2556 -482 -2554 1 a0_reg
rlabel metal1 -635 -2553 -633 -2551 3 a0
rlabel metal1 -742 -2561 -740 -2559 1 clk
rlabel metal1 -810 -2561 -809 -2559 1 clk
rlabel metal1 -829 -2510 -827 -2509 5 vdd
rlabel metal1 -835 -2582 -832 -2581 1 gnd
rlabel metal1 -833 -2561 -831 -2559 1 clk
rlabel metal1 -848 -2553 -846 -2551 3 b0
rlabel metal1 -698 -2556 -695 -2554 1 b0_reg
rlabel metal1 -605 -2890 -603 -2888 1 clk
rlabel metal1 -582 -2890 -581 -2888 1 clk
rlabel metal1 -514 -2890 -512 -2888 1 clk
rlabel metal1 -727 -2890 -725 -2888 1 clk
rlabel metal1 -795 -2890 -794 -2888 1 clk
rlabel metal1 -814 -2839 -812 -2838 5 vdd
rlabel metal1 -820 -2911 -817 -2910 1 gnd
rlabel metal1 -818 -2890 -816 -2888 1 clk
rlabel metal1 -581 -3157 -579 -3155 1 clk
rlabel metal1 -558 -3157 -557 -3155 1 clk
rlabel metal1 -490 -3157 -488 -3155 1 clk
rlabel metal1 -703 -3157 -701 -3155 1 clk
rlabel metal1 -771 -3157 -770 -3155 1 clk
rlabel metal1 -790 -3106 -788 -3105 5 vdd
rlabel metal1 -796 -3178 -793 -3177 1 gnd
rlabel metal1 -794 -3157 -792 -3155 1 clk
rlabel metal1 -765 -3467 -763 -3465 1 clk
rlabel metal1 -767 -3488 -764 -3487 1 gnd
rlabel metal1 -761 -3416 -759 -3415 5 vdd
rlabel metal1 -742 -3467 -741 -3465 1 clk
rlabel metal1 -674 -3467 -672 -3465 1 clk
rlabel metal1 -461 -3467 -459 -3465 1 clk
rlabel metal1 -529 -3467 -528 -3465 1 clk
rlabel metal1 -554 -3488 -551 -3487 1 gnd
rlabel metal1 -552 -3467 -550 -3465 1 clk
rlabel metal1 -620 -2882 -618 -2880 1 a1
rlabel metal1 -685 -2885 -680 -2883 1 b1_reg
rlabel metal1 -833 -2882 -831 -2880 1 b1
rlabel metal1 -470 -2885 -467 -2883 1 a1_reg
rlabel metal1 -62 -2891 -57 -2888 1 g1
rlabel metal1 -596 -3149 -594 -3147 1 a2
rlabel metal1 -446 -3152 -443 -3150 1 a2_reg
rlabel metal1 -659 -3152 -656 -3150 1 b2_reg
rlabel metal1 -809 -3149 -806 -3147 1 b2
rlabel metal1 -38 -3158 -33 -3155 1 g2
rlabel metal1 -9 -3468 -4 -3465 7 g3
rlabel metal1 -417 -3462 -414 -3460 1 a3_reg
rlabel metal1 -567 -3459 -564 -3457 1 a3
rlabel metal1 -630 -3462 -627 -3460 1 b3_reg
rlabel metal1 -780 -3459 -777 -3457 1 b3
rlabel metal1 200 -3519 203 -3516 1 help_c44
rlabel metal1 200 -3513 203 -3510 1 help_c43
rlabel metal1 198 -3432 201 -3429 1 help_c42
rlabel metal1 167 -3629 170 -3626 1 help_c44
rlabel metal1 106 -3628 109 -3625 1 p3
rlabel metal1 106 -3634 109 -3631 1 g2
rlabel metal1 160 -3599 160 -3599 5 vdd!
rlabel metal1 166 -3644 166 -3644 1 gnd!
rlabel metal1 130 -3657 130 -3657 1 gnd!
rlabel metal1 130 -3597 130 -3597 5 vdd!
rlabel metal1 194 -3174 197 -3171 1 help_c33
rlabel metal1 194 -3168 197 -3165 1 help_c32
rlabel metal1 192 -3081 195 -3078 1 help_c31
rlabel metal1 345 -2794 348 -2791 1 help_c21
rlabel metal1 407 -2789 410 -2786 7 c1
rlabel metal1 345 -2788 348 -2785 1 inter_c11
rlabel metal1 406 -2804 406 -2804 1 gnd!
rlabel metal1 400 -2759 400 -2759 5 vdd!
rlabel metal1 366 -2811 366 -2811 1 gnd!
rlabel metal1 363 -2746 363 -2746 5 vdd!
rlabel metal1 471 -3478 474 -3475 7 out_carry
rlabel metal1 409 -3483 412 -3480 1 help_c41
rlabel metal1 409 -3477 412 -3474 1 inter_c33
rlabel metal1 369 -3454 372 -3451 1 inter_c33
rlabel metal1 307 -3459 310 -3456 1 inter_c32
rlabel metal1 307 -3453 310 -3450 1 inter_c31
rlabel metal1 262 -3514 265 -3511 1 inter_c32
rlabel metal1 464 -3448 464 -3448 5 vdd!
rlabel metal1 427 -3435 427 -3435 5 vdd!
rlabel metal1 430 -3500 430 -3500 1 gnd!
rlabel metal1 470 -3493 470 -3493 1 gnd!
rlabel metal1 260 -3427 263 -3424 1 inter_c31
rlabel metal1 198 -3426 201 -3423 1 g3
rlabel metal1 167 -3547 170 -3544 1 help_c43
rlabel metal1 106 -3546 109 -3543 1 p3
rlabel metal1 106 -3552 109 -3549 1 help_c33
rlabel metal1 160 -3468 163 -3465 1 help_c42
rlabel metal1 99 -3473 102 -3470 1 p3
rlabel metal1 99 -3467 102 -3464 1 help_c32
rlabel metal1 96 -3351 99 -3348 1 p3
rlabel metal1 96 -3345 99 -3342 1 help_c31
rlabel metal1 157 -3346 160 -3343 1 help_c41
rlabel metal1 261 -3529 261 -3529 1 gnd!
rlabel metal1 221 -3536 221 -3536 1 gnd!
rlabel metal1 218 -3471 218 -3471 5 vdd!
rlabel metal1 120 -3314 120 -3314 5 vdd!
rlabel metal1 120 -3374 120 -3374 1 gnd!
rlabel metal1 150 -3316 150 -3316 5 vdd!
rlabel metal1 156 -3361 156 -3361 1 gnd!
rlabel metal1 123 -3436 123 -3436 5 vdd!
rlabel metal1 123 -3496 123 -3496 1 gnd!
rlabel metal1 159 -3483 159 -3483 1 gnd!
rlabel metal1 216 -3384 216 -3384 5 vdd!
rlabel metal1 219 -3449 219 -3449 1 gnd!
rlabel metal1 253 -3397 253 -3397 5 vdd!
rlabel metal1 259 -3442 259 -3442 1 gnd!
rlabel metal1 255 -3484 255 -3484 5 vdd!
rlabel metal1 153 -3438 153 -3438 5 vdd!
rlabel metal1 160 -3517 160 -3517 5 vdd!
rlabel metal1 166 -3562 166 -3562 1 gnd!
rlabel metal1 130 -3575 130 -3575 1 gnd!
rlabel metal1 130 -3515 130 -3515 5 vdd!
rlabel metal1 362 -3424 362 -3424 5 vdd!
rlabel metal1 325 -3411 325 -3411 5 vdd!
rlabel metal1 328 -3476 328 -3476 1 gnd!
rlabel metal1 368 -3469 368 -3469 1 gnd!
rlabel metal1 363 -3109 366 -3106 7 c2
rlabel metal1 301 -3108 304 -3105 1 inter_c21
rlabel metal1 301 -3114 304 -3111 1 inter_c22
rlabel metal1 256 -3169 259 -3166 1 inter_c22
rlabel metal1 254 -3082 257 -3079 1 inter_c21
rlabel metal1 192 -3087 195 -3084 1 g2
rlabel metal1 161 -3202 164 -3199 1 help_c33
rlabel metal1 100 -3207 103 -3204 1 g1
rlabel metal1 100 -3201 103 -3198 1 p2
rlabel metal1 154 -3123 157 -3120 1 help_c32
rlabel metal1 93 -3128 96 -3125 1 p2
rlabel metal1 93 -3122 96 -3119 1 help_c22
rlabel metal1 151 -3001 154 -2998 1 help_c31
rlabel metal1 90 -3006 93 -3003 1 p2
rlabel metal1 90 -3000 93 -2997 1 help_c21
rlabel metal1 362 -3124 362 -3124 1 gnd!
rlabel metal1 322 -3131 322 -3131 1 gnd!
rlabel metal1 319 -3066 319 -3066 5 vdd!
rlabel metal1 356 -3079 356 -3079 5 vdd!
rlabel metal1 124 -3170 124 -3170 5 vdd!
rlabel metal1 124 -3230 124 -3230 1 gnd!
rlabel metal1 160 -3217 160 -3217 1 gnd!
rlabel metal1 154 -3172 154 -3172 5 vdd!
rlabel metal1 147 -3093 147 -3093 5 vdd!
rlabel metal1 249 -3139 249 -3139 5 vdd!
rlabel metal1 253 -3097 253 -3097 1 gnd!
rlabel metal1 247 -3052 247 -3052 5 vdd!
rlabel metal1 213 -3104 213 -3104 1 gnd!
rlabel metal1 210 -3039 210 -3039 5 vdd!
rlabel metal1 153 -3138 153 -3138 1 gnd!
rlabel metal1 117 -3151 117 -3151 1 gnd!
rlabel metal1 117 -3091 117 -3091 5 vdd!
rlabel metal1 150 -3016 150 -3016 1 gnd!
rlabel metal1 144 -2971 144 -2971 5 vdd!
rlabel metal1 114 -3029 114 -3029 1 gnd!
rlabel metal1 114 -2969 114 -2969 5 vdd!
rlabel metal1 212 -3126 212 -3126 5 vdd!
rlabel metal1 215 -3191 215 -3191 1 gnd!
rlabel metal1 255 -3184 255 -3184 1 gnd!
rlabel metal1 256 -2818 259 -2815 7 inter_c11
rlabel metal1 194 -2817 197 -2814 1 help_c22
rlabel metal1 194 -2823 197 -2820 1 g1
rlabel metal1 156 -2859 159 -2856 1 help_c22
rlabel metal1 95 -2864 98 -2861 1 g0
rlabel metal1 95 -2858 98 -2855 1 p1
rlabel metal1 153 -2737 156 -2734 1 help_c21
rlabel metal1 92 -2736 95 -2733 1 p1
rlabel metal1 92 -2742 95 -2739 1 help_c1
rlabel metal1 116 -2705 116 -2705 5 vdd!
rlabel metal1 116 -2765 116 -2765 1 gnd!
rlabel metal1 146 -2707 146 -2707 5 vdd!
rlabel metal1 152 -2752 152 -2752 1 gnd!
rlabel metal1 119 -2827 119 -2827 5 vdd!
rlabel metal1 119 -2887 119 -2887 1 gnd!
rlabel metal1 149 -2829 149 -2829 5 vdd!
rlabel metal1 155 -2874 155 -2874 1 gnd!
rlabel metal1 212 -2775 212 -2775 5 vdd!
rlabel metal1 215 -2840 215 -2840 1 gnd!
rlabel metal1 249 -2788 249 -2788 5 vdd!
rlabel metal1 255 -2833 255 -2833 1 gnd!
rlabel metal1 109 -2462 109 -2462 5 vdd!
rlabel metal1 109 -2522 109 -2522 1 gnd!
rlabel metal1 139 -2464 139 -2464 5 vdd!
rlabel metal1 145 -2509 145 -2509 1 gnd!
rlabel metal1 202 -2410 202 -2410 5 vdd!
rlabel metal1 205 -2475 205 -2475 1 gnd!
rlabel metal1 239 -2423 239 -2423 5 vdd!
rlabel metal1 245 -2468 245 -2468 1 gnd!
rlabel metal1 85 -2499 88 -2496 3 p0
rlabel metal1 85 -2493 88 -2490 3 carry_reg
rlabel metal1 146 -2494 149 -2491 1 help_c1
rlabel metal1 184 -2458 187 -2455 1 g0
rlabel metal1 184 -2452 187 -2449 1 help_c1
rlabel metal1 246 -2453 249 -2450 7 c0
rlabel metal1 656 -2363 695 -2358 1 carry_reg
rlabel metal1 692 -3236 729 -3231 1 c2
rlabel metal1 686 -3315 702 -3309 1 p3
rlabel metal1 671 -2930 708 -2925 1 c1
rlabel metal1 665 -3009 681 -3003 1 p2
rlabel metal1 641 -2750 657 -2744 1 p1
rlabel metal1 647 -2671 684 -2666 1 c0
rlabel metal1 1006 -3278 1009 -3276 1 s3_reg
rlabel metal1 985 -2972 988 -2970 1 s2_reg
rlabel metal1 961 -2713 964 -2711 1 s1_reg
rlabel metal1 871 -3283 873 -3281 1 clk
rlabel metal1 869 -3304 872 -3303 1 gnd
rlabel metal1 875 -3232 877 -3231 5 vdd
rlabel metal1 894 -3283 895 -3281 1 clk
rlabel metal1 962 -3283 964 -3281 1 clk
rlabel metal1 604 -3217 718 -3212 5 VDD
rlabel metal1 580 -3379 694 -3373 1 GND
rlabel metal1 850 -2977 852 -2975 1 clk
rlabel metal1 848 -2998 851 -2997 1 gnd
rlabel metal1 854 -2926 856 -2925 5 vdd
rlabel metal1 873 -2977 874 -2975 1 clk
rlabel metal1 941 -2977 943 -2975 1 clk
rlabel metal1 583 -2911 697 -2906 5 VDD
rlabel metal1 559 -3073 673 -3067 1 GND
rlabel metal1 826 -2718 828 -2716 1 clk
rlabel metal1 824 -2739 827 -2738 1 gnd
rlabel metal1 830 -2667 832 -2666 5 vdd
rlabel metal1 849 -2718 850 -2716 1 clk
rlabel metal1 917 -2718 919 -2716 1 clk
rlabel metal1 559 -2652 673 -2647 5 VDD
rlabel metal1 535 -2814 649 -2808 1 GND
rlabel metal1 971 -2405 974 -2403 1 s0_reg
rlabel metal1 836 -2410 838 -2408 1 clk
rlabel metal1 834 -2431 837 -2430 1 gnd
rlabel metal1 840 -2359 842 -2358 5 vdd
rlabel metal1 859 -2410 860 -2408 1 clk
rlabel metal1 927 -2410 929 -2408 1 clk
rlabel metal1 651 -2442 667 -2436 1 p0
rlabel metal1 569 -2344 683 -2339 5 VDD
rlabel metal1 545 -2506 659 -2500 1 GND
rlabel metal1 65 -2347 68 -2345 1 carry_reg
rlabel metal1 -85 -2344 -83 -2342 1 carry
rlabel metal1 21 -2352 23 -2350 1 clk
rlabel metal1 -47 -2352 -46 -2350 1 clk
rlabel metal1 -66 -2301 -64 -2300 5 vdd
rlabel metal1 -72 -2373 -69 -2372 1 gnd
rlabel metal1 -70 -2352 -68 -2350 1 clk
rlabel metal1 611 -3485 613 -3483 1 clk
rlabel metal1 609 -3506 612 -3505 1 gnd
rlabel metal1 615 -3434 617 -3433 5 vdd
rlabel metal1 634 -3485 635 -3483 1 clk
rlabel metal1 702 -3485 704 -3483 1 clk
rlabel metal1 596 -3477 598 -3475 1 out_carry
rlabel metal1 745 -3480 750 -3478 1 out_carry_reg
rlabel metal1 -321 -2659 -315 -2654 1 p0
rlabel metal1 -306 -2986 -300 -2983 1 p1
rlabel metal1 -282 -3253 -276 -3250 1 p2
rlabel metal1 -253 -3564 -247 -3560 1 p3
<< end >>
