magic
tech scmos
timestamp 1732057525
<< nwell >>
rect -316 543 -282 579
rect -275 542 -251 566
rect -415 502 -381 526
rect -375 501 -351 525
rect -408 259 -374 283
rect -368 258 -344 282
rect -306 178 -272 214
rect -155 207 -121 243
rect -114 206 -90 230
rect -265 177 -241 201
rect -405 137 -371 161
rect -365 136 -341 160
rect -410 -5 -376 19
rect -370 -6 -346 18
rect -308 -86 -274 -50
rect -267 -87 -243 -63
rect -407 -127 -373 -103
rect -367 -128 -343 -104
rect -199 -113 -165 -77
rect -158 -114 -134 -90
rect -306 -173 -272 -137
rect -265 -174 -241 -150
rect -400 -206 -366 -182
rect -360 -207 -336 -183
rect -404 -350 -370 -326
rect -364 -351 -340 -327
rect -302 -431 -268 -395
rect -261 -432 -237 -408
rect -401 -472 -367 -448
rect -361 -473 -337 -449
rect -193 -458 -159 -422
rect -152 -459 -128 -435
rect -91 -482 -57 -446
rect -300 -518 -266 -482
rect -50 -483 -26 -459
rect -259 -519 -235 -495
rect -394 -551 -360 -527
rect -354 -552 -330 -528
rect -394 -633 -360 -609
rect -354 -634 -330 -610
<< ntransistor >>
rect -264 528 -262 534
rect -305 522 -303 528
rect -295 522 -293 528
rect -404 476 -402 488
rect -394 476 -392 488
rect -364 487 -362 493
rect -397 233 -395 245
rect -387 233 -385 245
rect -357 244 -355 250
rect -103 192 -101 198
rect -144 186 -142 192
rect -134 186 -132 192
rect -254 163 -252 169
rect -295 157 -293 163
rect -285 157 -283 163
rect -394 111 -392 123
rect -384 111 -382 123
rect -354 122 -352 128
rect -399 -31 -397 -19
rect -389 -31 -387 -19
rect -359 -20 -357 -14
rect -256 -101 -254 -95
rect -297 -107 -295 -101
rect -287 -107 -285 -101
rect -147 -128 -145 -122
rect -188 -134 -186 -128
rect -178 -134 -176 -128
rect -396 -153 -394 -141
rect -386 -153 -384 -141
rect -356 -142 -354 -136
rect -254 -188 -252 -182
rect -295 -194 -293 -188
rect -285 -194 -283 -188
rect -389 -232 -387 -220
rect -379 -232 -377 -220
rect -349 -221 -347 -215
rect -393 -376 -391 -364
rect -383 -376 -381 -364
rect -353 -365 -351 -359
rect -250 -446 -248 -440
rect -291 -452 -289 -446
rect -281 -452 -279 -446
rect -141 -473 -139 -467
rect -182 -479 -180 -473
rect -172 -479 -170 -473
rect -390 -498 -388 -486
rect -380 -498 -378 -486
rect -350 -487 -348 -481
rect -39 -497 -37 -491
rect -80 -503 -78 -497
rect -70 -503 -68 -497
rect -248 -533 -246 -527
rect -289 -539 -287 -533
rect -279 -539 -277 -533
rect -383 -577 -381 -565
rect -373 -577 -371 -565
rect -343 -566 -341 -560
rect -383 -659 -381 -647
rect -373 -659 -371 -647
rect -343 -648 -341 -642
<< ptransistor >>
rect -305 549 -303 573
rect -295 549 -293 573
rect -264 548 -262 560
rect -404 508 -402 520
rect -394 508 -392 520
rect -364 507 -362 519
rect -397 265 -395 277
rect -387 265 -385 277
rect -357 264 -355 276
rect -144 213 -142 237
rect -134 213 -132 237
rect -295 184 -293 208
rect -285 184 -283 208
rect -254 183 -252 195
rect -103 212 -101 224
rect -394 143 -392 155
rect -384 143 -382 155
rect -354 142 -352 154
rect -399 1 -397 13
rect -389 1 -387 13
rect -359 0 -357 12
rect -297 -80 -295 -56
rect -287 -80 -285 -56
rect -256 -81 -254 -69
rect -188 -107 -186 -83
rect -178 -107 -176 -83
rect -396 -121 -394 -109
rect -386 -121 -384 -109
rect -356 -122 -354 -110
rect -147 -108 -145 -96
rect -295 -167 -293 -143
rect -285 -167 -283 -143
rect -389 -200 -387 -188
rect -379 -200 -377 -188
rect -254 -168 -252 -156
rect -349 -201 -347 -189
rect -393 -344 -391 -332
rect -383 -344 -381 -332
rect -353 -345 -351 -333
rect -291 -425 -289 -401
rect -281 -425 -279 -401
rect -250 -426 -248 -414
rect -182 -452 -180 -428
rect -172 -452 -170 -428
rect -390 -466 -388 -454
rect -380 -466 -378 -454
rect -350 -467 -348 -455
rect -141 -453 -139 -441
rect -80 -476 -78 -452
rect -70 -476 -68 -452
rect -289 -512 -287 -488
rect -279 -512 -277 -488
rect -39 -477 -37 -465
rect -383 -545 -381 -533
rect -373 -545 -371 -533
rect -248 -513 -246 -501
rect -343 -546 -341 -534
rect -383 -627 -381 -615
rect -373 -627 -371 -615
rect -343 -628 -341 -616
<< ndiffusion >>
rect -265 528 -264 534
rect -262 528 -261 534
rect -306 522 -305 528
rect -303 522 -301 528
rect -297 522 -295 528
rect -293 522 -292 528
rect -405 476 -404 488
rect -402 476 -394 488
rect -392 476 -391 488
rect -365 487 -364 493
rect -362 487 -361 493
rect -398 233 -397 245
rect -395 233 -387 245
rect -385 233 -384 245
rect -358 244 -357 250
rect -355 244 -354 250
rect -104 192 -103 198
rect -101 192 -100 198
rect -145 186 -144 192
rect -142 186 -140 192
rect -136 186 -134 192
rect -132 186 -131 192
rect -255 163 -254 169
rect -252 163 -251 169
rect -296 157 -295 163
rect -293 157 -291 163
rect -287 157 -285 163
rect -283 157 -282 163
rect -395 111 -394 123
rect -392 111 -384 123
rect -382 111 -381 123
rect -355 122 -354 128
rect -352 122 -351 128
rect -400 -31 -399 -19
rect -397 -31 -389 -19
rect -387 -31 -386 -19
rect -360 -20 -359 -14
rect -357 -20 -356 -14
rect -257 -101 -256 -95
rect -254 -101 -253 -95
rect -298 -107 -297 -101
rect -295 -107 -293 -101
rect -289 -107 -287 -101
rect -285 -107 -284 -101
rect -148 -128 -147 -122
rect -145 -128 -144 -122
rect -189 -134 -188 -128
rect -186 -134 -184 -128
rect -180 -134 -178 -128
rect -176 -134 -175 -128
rect -397 -153 -396 -141
rect -394 -153 -386 -141
rect -384 -153 -383 -141
rect -357 -142 -356 -136
rect -354 -142 -353 -136
rect -255 -188 -254 -182
rect -252 -188 -251 -182
rect -296 -194 -295 -188
rect -293 -194 -291 -188
rect -287 -194 -285 -188
rect -283 -194 -282 -188
rect -390 -232 -389 -220
rect -387 -232 -379 -220
rect -377 -232 -376 -220
rect -350 -221 -349 -215
rect -347 -221 -346 -215
rect -394 -376 -393 -364
rect -391 -376 -383 -364
rect -381 -376 -380 -364
rect -354 -365 -353 -359
rect -351 -365 -350 -359
rect -251 -446 -250 -440
rect -248 -446 -247 -440
rect -292 -452 -291 -446
rect -289 -452 -287 -446
rect -283 -452 -281 -446
rect -279 -452 -278 -446
rect -142 -473 -141 -467
rect -139 -473 -138 -467
rect -183 -479 -182 -473
rect -180 -479 -178 -473
rect -174 -479 -172 -473
rect -170 -479 -169 -473
rect -391 -498 -390 -486
rect -388 -498 -380 -486
rect -378 -498 -377 -486
rect -351 -487 -350 -481
rect -348 -487 -347 -481
rect -40 -497 -39 -491
rect -37 -497 -36 -491
rect -81 -503 -80 -497
rect -78 -503 -76 -497
rect -72 -503 -70 -497
rect -68 -503 -67 -497
rect -249 -533 -248 -527
rect -246 -533 -245 -527
rect -290 -539 -289 -533
rect -287 -539 -285 -533
rect -281 -539 -279 -533
rect -277 -539 -276 -533
rect -384 -577 -383 -565
rect -381 -577 -373 -565
rect -371 -577 -370 -565
rect -344 -566 -343 -560
rect -341 -566 -340 -560
rect -384 -659 -383 -647
rect -381 -659 -373 -647
rect -371 -659 -370 -647
rect -344 -648 -343 -642
rect -341 -648 -340 -642
<< pdiffusion >>
rect -306 549 -305 573
rect -303 549 -295 573
rect -293 549 -292 573
rect -265 548 -264 560
rect -262 548 -261 560
rect -405 508 -404 520
rect -402 508 -400 520
rect -396 508 -394 520
rect -392 508 -391 520
rect -365 507 -364 519
rect -362 507 -361 519
rect -398 265 -397 277
rect -395 265 -393 277
rect -389 265 -387 277
rect -385 265 -384 277
rect -358 264 -357 276
rect -355 264 -354 276
rect -145 213 -144 237
rect -142 213 -134 237
rect -132 213 -131 237
rect -296 184 -295 208
rect -293 184 -285 208
rect -283 184 -282 208
rect -255 183 -254 195
rect -252 183 -251 195
rect -104 212 -103 224
rect -101 212 -100 224
rect -395 143 -394 155
rect -392 143 -390 155
rect -386 143 -384 155
rect -382 143 -381 155
rect -355 142 -354 154
rect -352 142 -351 154
rect -400 1 -399 13
rect -397 1 -395 13
rect -391 1 -389 13
rect -387 1 -386 13
rect -360 0 -359 12
rect -357 0 -356 12
rect -298 -80 -297 -56
rect -295 -80 -287 -56
rect -285 -80 -284 -56
rect -257 -81 -256 -69
rect -254 -81 -253 -69
rect -189 -107 -188 -83
rect -186 -107 -178 -83
rect -176 -107 -175 -83
rect -397 -121 -396 -109
rect -394 -121 -392 -109
rect -388 -121 -386 -109
rect -384 -121 -383 -109
rect -357 -122 -356 -110
rect -354 -122 -353 -110
rect -148 -108 -147 -96
rect -145 -108 -144 -96
rect -296 -167 -295 -143
rect -293 -167 -285 -143
rect -283 -167 -282 -143
rect -390 -200 -389 -188
rect -387 -200 -385 -188
rect -381 -200 -379 -188
rect -377 -200 -376 -188
rect -255 -168 -254 -156
rect -252 -168 -251 -156
rect -350 -201 -349 -189
rect -347 -201 -346 -189
rect -394 -344 -393 -332
rect -391 -344 -389 -332
rect -385 -344 -383 -332
rect -381 -344 -380 -332
rect -354 -345 -353 -333
rect -351 -345 -350 -333
rect -292 -425 -291 -401
rect -289 -425 -281 -401
rect -279 -425 -278 -401
rect -251 -426 -250 -414
rect -248 -426 -247 -414
rect -183 -452 -182 -428
rect -180 -452 -172 -428
rect -170 -452 -169 -428
rect -391 -466 -390 -454
rect -388 -466 -386 -454
rect -382 -466 -380 -454
rect -378 -466 -377 -454
rect -351 -467 -350 -455
rect -348 -467 -347 -455
rect -142 -453 -141 -441
rect -139 -453 -138 -441
rect -81 -476 -80 -452
rect -78 -476 -70 -452
rect -68 -476 -67 -452
rect -290 -512 -289 -488
rect -287 -512 -279 -488
rect -277 -512 -276 -488
rect -40 -477 -39 -465
rect -37 -477 -36 -465
rect -384 -545 -383 -533
rect -381 -545 -379 -533
rect -375 -545 -373 -533
rect -371 -545 -370 -533
rect -249 -513 -248 -501
rect -246 -513 -245 -501
rect -344 -546 -343 -534
rect -341 -546 -340 -534
rect -384 -627 -383 -615
rect -381 -627 -379 -615
rect -375 -627 -373 -615
rect -371 -627 -370 -615
rect -344 -628 -343 -616
rect -341 -628 -340 -616
<< ndcontact >>
rect -269 528 -265 534
rect -261 528 -257 534
rect -310 522 -306 528
rect -301 522 -297 528
rect -292 522 -288 528
rect -409 476 -405 488
rect -391 476 -387 488
rect -369 487 -365 493
rect -361 487 -357 493
rect -402 233 -398 245
rect -384 233 -380 245
rect -362 244 -358 250
rect -354 244 -350 250
rect -108 192 -104 198
rect -100 192 -96 198
rect -149 186 -145 192
rect -140 186 -136 192
rect -131 186 -127 192
rect -259 163 -255 169
rect -251 163 -247 169
rect -300 157 -296 163
rect -291 157 -287 163
rect -282 157 -278 163
rect -399 111 -395 123
rect -381 111 -377 123
rect -359 122 -355 128
rect -351 122 -347 128
rect -404 -31 -400 -19
rect -386 -31 -382 -19
rect -364 -20 -360 -14
rect -356 -20 -352 -14
rect -261 -101 -257 -95
rect -253 -101 -249 -95
rect -302 -107 -298 -101
rect -293 -107 -289 -101
rect -284 -107 -280 -101
rect -152 -128 -148 -122
rect -144 -128 -140 -122
rect -193 -134 -189 -128
rect -184 -134 -180 -128
rect -175 -134 -171 -128
rect -401 -153 -397 -141
rect -383 -153 -379 -141
rect -361 -142 -357 -136
rect -353 -142 -349 -136
rect -259 -188 -255 -182
rect -251 -188 -247 -182
rect -300 -194 -296 -188
rect -291 -194 -287 -188
rect -282 -194 -278 -188
rect -394 -232 -390 -220
rect -376 -232 -372 -220
rect -354 -221 -350 -215
rect -346 -221 -342 -215
rect -398 -376 -394 -364
rect -380 -376 -376 -364
rect -358 -365 -354 -359
rect -350 -365 -346 -359
rect -255 -446 -251 -440
rect -247 -446 -243 -440
rect -296 -452 -292 -446
rect -287 -452 -283 -446
rect -278 -452 -274 -446
rect -146 -473 -142 -467
rect -138 -473 -134 -467
rect -187 -479 -183 -473
rect -178 -479 -174 -473
rect -169 -479 -165 -473
rect -395 -498 -391 -486
rect -377 -498 -373 -486
rect -355 -487 -351 -481
rect -347 -487 -343 -481
rect -44 -497 -40 -491
rect -36 -497 -32 -491
rect -85 -503 -81 -497
rect -76 -503 -72 -497
rect -67 -503 -63 -497
rect -253 -533 -249 -527
rect -245 -533 -241 -527
rect -294 -539 -290 -533
rect -285 -539 -281 -533
rect -276 -539 -272 -533
rect -388 -577 -384 -565
rect -370 -577 -366 -565
rect -348 -566 -344 -560
rect -340 -566 -336 -560
rect -388 -659 -384 -647
rect -370 -659 -366 -647
rect -348 -648 -344 -642
rect -340 -648 -336 -642
<< pdcontact >>
rect -310 549 -306 573
rect -292 549 -288 573
rect -269 548 -265 560
rect -261 548 -257 560
rect -409 508 -405 520
rect -400 508 -396 520
rect -391 508 -387 520
rect -369 507 -365 519
rect -361 507 -357 519
rect -402 265 -398 277
rect -393 265 -389 277
rect -384 265 -380 277
rect -362 264 -358 276
rect -354 264 -350 276
rect -149 213 -145 237
rect -131 213 -127 237
rect -300 184 -296 208
rect -282 184 -278 208
rect -259 183 -255 195
rect -251 183 -247 195
rect -108 212 -104 224
rect -100 212 -96 224
rect -399 143 -395 155
rect -390 143 -386 155
rect -381 143 -377 155
rect -359 142 -355 154
rect -351 142 -347 154
rect -404 1 -400 13
rect -395 1 -391 13
rect -386 1 -382 13
rect -364 0 -360 12
rect -356 0 -352 12
rect -302 -80 -298 -56
rect -284 -80 -280 -56
rect -261 -81 -257 -69
rect -253 -81 -249 -69
rect -193 -107 -189 -83
rect -175 -107 -171 -83
rect -401 -121 -397 -109
rect -392 -121 -388 -109
rect -383 -121 -379 -109
rect -361 -122 -357 -110
rect -353 -122 -349 -110
rect -152 -108 -148 -96
rect -144 -108 -140 -96
rect -300 -167 -296 -143
rect -282 -167 -278 -143
rect -394 -200 -390 -188
rect -385 -200 -381 -188
rect -376 -200 -372 -188
rect -259 -168 -255 -156
rect -251 -168 -247 -156
rect -354 -201 -350 -189
rect -346 -201 -342 -189
rect -398 -344 -394 -332
rect -389 -344 -385 -332
rect -380 -344 -376 -332
rect -358 -345 -354 -333
rect -350 -345 -346 -333
rect -296 -425 -292 -401
rect -278 -425 -274 -401
rect -255 -426 -251 -414
rect -247 -426 -243 -414
rect -187 -452 -183 -428
rect -169 -452 -165 -428
rect -395 -466 -391 -454
rect -386 -466 -382 -454
rect -377 -466 -373 -454
rect -355 -467 -351 -455
rect -347 -467 -343 -455
rect -146 -453 -142 -441
rect -138 -453 -134 -441
rect -85 -476 -81 -452
rect -67 -476 -63 -452
rect -294 -512 -290 -488
rect -276 -512 -272 -488
rect -44 -477 -40 -465
rect -36 -477 -32 -465
rect -388 -545 -384 -533
rect -379 -545 -375 -533
rect -370 -545 -366 -533
rect -253 -513 -249 -501
rect -245 -513 -241 -501
rect -348 -546 -344 -534
rect -340 -546 -336 -534
rect -388 -627 -384 -615
rect -379 -627 -375 -615
rect -370 -627 -366 -615
rect -348 -628 -344 -616
rect -340 -628 -336 -616
<< polysilicon >>
rect -305 573 -303 576
rect -295 573 -293 576
rect -264 560 -262 563
rect -305 528 -303 549
rect -295 528 -293 549
rect -264 534 -262 548
rect -404 520 -402 523
rect -394 520 -392 523
rect -264 525 -262 528
rect -364 519 -362 522
rect -305 519 -303 522
rect -295 519 -293 522
rect -404 488 -402 508
rect -394 488 -392 508
rect -364 493 -362 507
rect -364 484 -362 487
rect -404 473 -402 476
rect -394 473 -392 476
rect -397 277 -395 280
rect -387 277 -385 280
rect -357 276 -355 279
rect -397 245 -395 265
rect -387 245 -385 265
rect -357 250 -355 264
rect -357 241 -355 244
rect -144 237 -142 240
rect -134 237 -132 240
rect -397 230 -395 233
rect -387 230 -385 233
rect -103 224 -101 227
rect -295 208 -293 211
rect -285 208 -283 211
rect -254 195 -252 198
rect -295 163 -293 184
rect -285 163 -283 184
rect -144 192 -142 213
rect -134 192 -132 213
rect -103 198 -101 212
rect -103 189 -101 192
rect -144 183 -142 186
rect -134 183 -132 186
rect -254 169 -252 183
rect -394 155 -392 158
rect -384 155 -382 158
rect -254 160 -252 163
rect -354 154 -352 157
rect -295 154 -293 157
rect -285 154 -283 157
rect -394 123 -392 143
rect -384 123 -382 143
rect -354 128 -352 142
rect -354 119 -352 122
rect -394 108 -392 111
rect -384 108 -382 111
rect -399 13 -397 16
rect -389 13 -387 16
rect -359 12 -357 15
rect -399 -19 -397 1
rect -389 -19 -387 1
rect -359 -14 -357 0
rect -359 -23 -357 -20
rect -399 -34 -397 -31
rect -389 -34 -387 -31
rect -297 -56 -295 -53
rect -287 -56 -285 -53
rect -256 -69 -254 -66
rect -297 -101 -295 -80
rect -287 -101 -285 -80
rect -256 -95 -254 -81
rect -188 -83 -186 -80
rect -178 -83 -176 -80
rect -396 -109 -394 -106
rect -386 -109 -384 -106
rect -256 -104 -254 -101
rect -147 -96 -145 -93
rect -356 -110 -354 -107
rect -297 -110 -295 -107
rect -287 -110 -285 -107
rect -396 -141 -394 -121
rect -386 -141 -384 -121
rect -356 -136 -354 -122
rect -188 -128 -186 -107
rect -178 -128 -176 -107
rect -147 -122 -145 -108
rect -147 -131 -145 -128
rect -188 -137 -186 -134
rect -178 -137 -176 -134
rect -356 -145 -354 -142
rect -295 -143 -293 -140
rect -285 -143 -283 -140
rect -396 -156 -394 -153
rect -386 -156 -384 -153
rect -254 -156 -252 -153
rect -389 -188 -387 -185
rect -379 -188 -377 -185
rect -349 -189 -347 -186
rect -295 -188 -293 -167
rect -285 -188 -283 -167
rect -254 -182 -252 -168
rect -389 -220 -387 -200
rect -379 -220 -377 -200
rect -254 -191 -252 -188
rect -295 -197 -293 -194
rect -285 -197 -283 -194
rect -349 -215 -347 -201
rect -349 -224 -347 -221
rect -389 -235 -387 -232
rect -379 -235 -377 -232
rect -393 -332 -391 -329
rect -383 -332 -381 -329
rect -353 -333 -351 -330
rect -393 -364 -391 -344
rect -383 -364 -381 -344
rect -353 -359 -351 -345
rect -353 -368 -351 -365
rect -393 -379 -391 -376
rect -383 -379 -381 -376
rect -291 -401 -289 -398
rect -281 -401 -279 -398
rect -250 -414 -248 -411
rect -291 -446 -289 -425
rect -281 -446 -279 -425
rect -250 -440 -248 -426
rect -182 -428 -180 -425
rect -172 -428 -170 -425
rect -390 -454 -388 -451
rect -380 -454 -378 -451
rect -250 -449 -248 -446
rect -141 -441 -139 -438
rect -350 -455 -348 -452
rect -291 -455 -289 -452
rect -281 -455 -279 -452
rect -390 -486 -388 -466
rect -380 -486 -378 -466
rect -350 -481 -348 -467
rect -182 -473 -180 -452
rect -172 -473 -170 -452
rect -80 -452 -78 -449
rect -70 -452 -68 -449
rect -141 -467 -139 -453
rect -141 -476 -139 -473
rect -39 -465 -37 -462
rect -182 -482 -180 -479
rect -172 -482 -170 -479
rect -350 -490 -348 -487
rect -289 -488 -287 -485
rect -279 -488 -277 -485
rect -390 -501 -388 -498
rect -380 -501 -378 -498
rect -80 -497 -78 -476
rect -70 -497 -68 -476
rect -39 -491 -37 -477
rect -248 -501 -246 -498
rect -383 -533 -381 -530
rect -373 -533 -371 -530
rect -343 -534 -341 -531
rect -289 -533 -287 -512
rect -279 -533 -277 -512
rect -39 -500 -37 -497
rect -80 -506 -78 -503
rect -70 -506 -68 -503
rect -248 -527 -246 -513
rect -383 -565 -381 -545
rect -373 -565 -371 -545
rect -248 -536 -246 -533
rect -289 -542 -287 -539
rect -279 -542 -277 -539
rect -343 -560 -341 -546
rect -343 -569 -341 -566
rect -383 -580 -381 -577
rect -373 -580 -371 -577
rect -383 -615 -381 -612
rect -373 -615 -371 -612
rect -343 -616 -341 -613
rect -383 -647 -381 -627
rect -373 -647 -371 -627
rect -343 -642 -341 -628
rect -343 -651 -341 -648
rect -383 -662 -381 -659
rect -373 -662 -371 -659
<< polycontact >>
rect -309 531 -305 535
rect -299 538 -295 542
rect -268 537 -264 541
rect -408 497 -404 501
rect -398 491 -394 495
rect -368 496 -364 500
rect -401 254 -397 258
rect -391 248 -387 252
rect -361 253 -357 257
rect -148 195 -144 199
rect -299 166 -295 170
rect -289 173 -285 177
rect -138 202 -134 206
rect -107 201 -103 205
rect -258 172 -254 176
rect -398 132 -394 136
rect -388 126 -384 130
rect -358 131 -354 135
rect -403 -10 -399 -6
rect -393 -16 -389 -12
rect -363 -11 -359 -7
rect -301 -98 -297 -94
rect -291 -91 -287 -87
rect -260 -92 -256 -88
rect -400 -132 -396 -128
rect -390 -138 -386 -134
rect -360 -133 -356 -129
rect -192 -125 -188 -121
rect -182 -118 -178 -114
rect -151 -119 -147 -115
rect -299 -185 -295 -181
rect -289 -178 -285 -174
rect -258 -179 -254 -175
rect -393 -211 -389 -207
rect -383 -217 -379 -213
rect -353 -212 -349 -208
rect -397 -355 -393 -351
rect -387 -361 -383 -357
rect -357 -356 -353 -352
rect -295 -443 -291 -439
rect -285 -436 -281 -432
rect -254 -437 -250 -433
rect -394 -477 -390 -473
rect -384 -483 -380 -479
rect -354 -478 -350 -474
rect -186 -470 -182 -466
rect -176 -463 -172 -459
rect -145 -464 -141 -460
rect -84 -494 -80 -490
rect -74 -487 -70 -483
rect -43 -488 -39 -484
rect -293 -530 -289 -526
rect -283 -523 -279 -519
rect -252 -524 -248 -520
rect -387 -556 -383 -552
rect -377 -562 -373 -558
rect -347 -557 -343 -553
rect -387 -638 -383 -634
rect -377 -644 -373 -640
rect -347 -639 -343 -635
<< metal1 >>
rect -354 579 -274 582
rect -415 528 -372 529
rect -354 528 -351 579
rect -310 573 -307 579
rect -277 569 -274 579
rect -277 566 -251 569
rect -415 526 -351 528
rect -409 520 -406 526
rect -390 520 -387 526
rect -375 525 -351 526
rect -334 538 -299 541
rect -291 540 -288 549
rect -269 560 -266 566
rect -369 519 -366 525
rect -400 505 -397 508
rect -400 502 -387 505
rect -415 497 -408 500
rect -390 499 -387 502
rect -390 496 -368 499
rect -360 499 -357 507
rect -334 499 -329 538
rect -291 537 -268 540
rect -260 540 -257 548
rect -260 537 -251 540
rect -316 532 -309 535
rect -291 534 -288 537
rect -260 534 -257 537
rect -300 531 -288 534
rect -300 528 -297 531
rect -269 524 -266 528
rect -310 516 -307 522
rect -291 516 -288 522
rect -279 521 -251 524
rect -279 516 -275 521
rect -360 496 -329 499
rect -318 513 -275 516
rect -415 491 -398 494
rect -390 488 -387 496
rect -360 493 -357 496
rect -369 483 -366 487
rect -318 483 -314 513
rect -379 480 -314 483
rect -409 470 -406 476
rect -379 470 -375 480
rect -415 467 -375 470
rect -408 285 -365 286
rect -345 285 -302 286
rect -408 283 -302 285
rect -402 277 -399 283
rect -383 277 -380 283
rect -368 282 -302 283
rect -362 276 -359 282
rect -393 262 -390 265
rect -393 259 -380 262
rect -408 254 -401 257
rect -383 256 -380 259
rect -383 253 -361 256
rect -353 256 -350 264
rect -353 253 -333 256
rect -434 248 -391 251
rect -383 245 -380 253
rect -353 250 -350 253
rect -362 240 -359 244
rect -372 237 -344 240
rect -402 227 -399 233
rect -372 227 -368 237
rect -408 224 -368 227
rect -306 217 -302 282
rect -243 246 -154 247
rect -243 243 -113 246
rect -306 214 -264 217
rect -300 208 -297 214
rect -267 204 -264 214
rect -243 205 -240 243
rect -149 237 -146 243
rect -116 233 -113 243
rect -116 230 -90 233
rect -244 204 -240 205
rect -267 202 -240 204
rect -205 202 -138 205
rect -130 204 -127 213
rect -108 224 -105 230
rect -267 201 -241 202
rect -325 173 -289 176
rect -281 175 -278 184
rect -259 195 -256 201
rect -405 163 -362 164
rect -405 161 -341 163
rect -399 155 -396 161
rect -380 155 -377 161
rect -365 160 -341 161
rect -359 154 -356 160
rect -390 140 -387 143
rect -390 137 -377 140
rect -405 132 -398 135
rect -380 134 -377 137
rect -380 131 -358 134
rect -350 134 -347 142
rect -325 134 -322 173
rect -281 172 -258 175
rect -250 175 -247 183
rect -205 175 -201 202
rect -130 201 -107 204
rect -99 204 -96 212
rect -99 201 -90 204
rect -170 196 -148 199
rect -130 198 -127 201
rect -99 198 -96 201
rect -139 195 -127 198
rect -139 192 -136 195
rect -108 188 -105 192
rect -149 180 -146 186
rect -130 180 -127 186
rect -118 185 -90 188
rect -118 180 -114 185
rect -250 172 -201 175
rect -161 177 -114 180
rect -306 167 -299 170
rect -281 169 -278 172
rect -250 169 -247 172
rect -290 166 -278 169
rect -290 163 -287 166
rect -259 159 -256 163
rect -161 159 -158 177
rect -300 151 -297 157
rect -281 151 -278 157
rect -269 156 -178 159
rect -175 156 -158 159
rect -269 151 -265 156
rect -350 131 -322 134
rect -310 148 -265 151
rect -405 126 -388 129
rect -380 123 -377 131
rect -350 128 -347 131
rect -359 118 -356 122
rect -310 118 -306 148
rect -369 115 -306 118
rect -399 105 -396 111
rect -369 105 -365 115
rect -405 102 -365 105
rect -410 21 -367 22
rect -410 19 -346 21
rect -404 13 -401 19
rect -385 13 -382 19
rect -370 18 -346 19
rect -364 12 -361 18
rect -395 -2 -392 1
rect -395 -5 -382 -2
rect -448 -10 -403 -7
rect -385 -8 -382 -5
rect -385 -11 -363 -8
rect -355 -8 -352 0
rect -355 -11 -335 -8
rect -410 -16 -393 -13
rect -385 -19 -382 -11
rect -355 -14 -352 -11
rect -364 -24 -361 -20
rect -374 -27 -346 -24
rect -404 -37 -401 -31
rect -374 -37 -370 -27
rect -410 -40 -370 -37
rect -338 -88 -335 -11
rect -308 -50 -266 -47
rect -302 -56 -299 -50
rect -269 -60 -266 -50
rect -269 -63 -243 -60
rect -338 -91 -291 -88
rect -283 -89 -280 -80
rect -261 -69 -258 -63
rect -199 -77 -157 -74
rect -283 -92 -260 -89
rect -252 -89 -249 -81
rect -193 -83 -190 -77
rect -252 -92 -230 -89
rect -308 -97 -301 -94
rect -283 -95 -280 -92
rect -252 -95 -249 -92
rect -292 -98 -280 -95
rect -407 -101 -364 -100
rect -292 -101 -289 -98
rect -407 -103 -343 -101
rect -401 -109 -398 -103
rect -382 -109 -379 -103
rect -367 -104 -343 -103
rect -361 -110 -358 -104
rect -261 -105 -258 -101
rect -392 -124 -389 -121
rect -302 -113 -299 -107
rect -283 -113 -280 -107
rect -271 -108 -243 -105
rect -271 -113 -267 -108
rect -308 -116 -267 -113
rect -233 -115 -230 -92
rect -160 -87 -157 -77
rect -160 -90 -134 -87
rect -233 -118 -182 -115
rect -174 -116 -171 -107
rect -152 -96 -149 -90
rect -174 -119 -151 -116
rect -143 -116 -140 -108
rect -143 -119 -134 -116
rect -392 -127 -379 -124
rect -483 -129 -477 -127
rect -483 -132 -400 -129
rect -382 -130 -379 -127
rect -382 -133 -360 -130
rect -352 -130 -349 -122
rect -236 -124 -192 -121
rect -352 -133 -332 -130
rect -407 -138 -390 -135
rect -382 -141 -379 -133
rect -352 -136 -349 -133
rect -361 -146 -358 -142
rect -371 -149 -343 -146
rect -401 -159 -398 -153
rect -371 -159 -367 -149
rect -407 -162 -367 -159
rect -335 -174 -332 -133
rect -306 -137 -264 -134
rect -300 -143 -297 -137
rect -267 -147 -264 -137
rect -267 -150 -241 -147
rect -335 -175 -330 -174
rect -335 -177 -289 -175
rect -333 -178 -289 -177
rect -281 -176 -278 -167
rect -259 -156 -256 -150
rect -281 -179 -258 -176
rect -250 -176 -247 -168
rect -236 -176 -233 -124
rect -174 -122 -171 -119
rect -143 -122 -140 -119
rect -183 -125 -171 -122
rect -183 -128 -180 -125
rect -152 -132 -149 -128
rect -193 -140 -190 -134
rect -174 -140 -171 -134
rect -162 -135 -134 -132
rect -162 -140 -158 -135
rect -199 -143 -158 -140
rect -250 -179 -233 -176
rect -400 -180 -357 -179
rect -400 -182 -336 -180
rect -394 -188 -391 -182
rect -375 -188 -372 -182
rect -360 -183 -336 -182
rect -354 -189 -351 -183
rect -319 -184 -299 -181
rect -385 -203 -382 -200
rect -385 -206 -372 -203
rect -400 -211 -393 -208
rect -375 -209 -372 -206
rect -375 -212 -353 -209
rect -345 -209 -342 -201
rect -319 -209 -315 -184
rect -281 -182 -278 -179
rect -250 -182 -247 -179
rect -290 -185 -278 -182
rect -290 -188 -287 -185
rect -259 -192 -256 -188
rect -300 -200 -297 -194
rect -281 -200 -278 -194
rect -269 -195 -241 -192
rect -269 -200 -265 -195
rect -306 -203 -265 -200
rect -345 -212 -315 -209
rect -400 -217 -383 -214
rect -375 -220 -372 -212
rect -345 -215 -342 -212
rect -354 -225 -351 -221
rect -364 -228 -336 -225
rect -394 -238 -391 -232
rect -364 -238 -360 -228
rect -400 -241 -360 -238
rect -404 -324 -361 -323
rect -404 -326 -340 -324
rect -398 -332 -395 -326
rect -379 -332 -376 -326
rect -364 -327 -340 -326
rect -358 -333 -355 -327
rect -389 -347 -386 -344
rect -389 -350 -376 -347
rect -456 -355 -397 -352
rect -379 -353 -376 -350
rect -379 -356 -357 -353
rect -349 -353 -346 -345
rect -349 -356 -96 -353
rect -404 -361 -387 -358
rect -379 -364 -376 -356
rect -349 -359 -346 -356
rect -270 -357 -96 -356
rect -104 -363 -96 -357
rect -358 -369 -355 -365
rect -368 -372 -340 -369
rect -398 -382 -395 -376
rect -368 -382 -364 -372
rect -404 -385 -364 -382
rect -302 -395 -260 -392
rect -296 -401 -293 -395
rect -263 -405 -260 -395
rect -263 -408 -237 -405
rect -302 -436 -285 -433
rect -277 -434 -274 -425
rect -255 -414 -252 -408
rect -193 -422 -151 -419
rect -277 -437 -254 -434
rect -246 -434 -243 -426
rect -187 -428 -184 -422
rect -246 -437 -225 -434
rect -314 -442 -295 -439
rect -401 -446 -358 -445
rect -401 -448 -337 -446
rect -395 -454 -392 -448
rect -376 -454 -373 -448
rect -361 -449 -337 -448
rect -355 -455 -352 -449
rect -386 -469 -383 -466
rect -386 -472 -373 -469
rect -444 -477 -394 -474
rect -376 -475 -373 -472
rect -376 -478 -354 -475
rect -346 -475 -343 -467
rect -314 -475 -311 -442
rect -277 -440 -274 -437
rect -246 -440 -243 -437
rect -286 -443 -274 -440
rect -286 -446 -283 -443
rect -255 -450 -252 -446
rect -296 -458 -293 -452
rect -277 -458 -274 -452
rect -265 -453 -237 -450
rect -265 -458 -261 -453
rect -302 -461 -261 -458
rect -229 -460 -225 -437
rect -154 -432 -151 -422
rect -154 -435 -128 -432
rect -229 -463 -176 -460
rect -168 -461 -165 -452
rect -146 -441 -143 -435
rect -91 -446 -49 -443
rect -168 -464 -145 -461
rect -137 -461 -134 -453
rect -85 -452 -82 -446
rect -137 -464 -119 -461
rect -346 -478 -311 -475
rect -206 -469 -186 -466
rect -401 -483 -384 -480
rect -376 -486 -373 -478
rect -346 -481 -343 -478
rect -300 -482 -258 -479
rect -355 -491 -352 -487
rect -294 -488 -291 -482
rect -365 -494 -337 -491
rect -395 -504 -392 -498
rect -365 -504 -361 -494
rect -401 -507 -361 -504
rect -261 -492 -258 -482
rect -261 -495 -235 -492
rect -326 -523 -283 -520
rect -275 -521 -272 -512
rect -253 -501 -250 -495
rect -394 -525 -351 -524
rect -394 -527 -330 -525
rect -388 -533 -385 -527
rect -369 -533 -366 -527
rect -354 -528 -330 -527
rect -348 -534 -345 -528
rect -379 -548 -376 -545
rect -379 -551 -366 -548
rect -394 -556 -387 -553
rect -369 -554 -366 -551
rect -369 -557 -347 -554
rect -339 -554 -336 -546
rect -326 -554 -323 -523
rect -275 -524 -252 -521
rect -244 -521 -241 -513
rect -206 -521 -202 -469
rect -168 -467 -165 -464
rect -137 -467 -134 -464
rect -177 -470 -165 -467
rect -177 -473 -174 -470
rect -146 -477 -143 -473
rect -187 -485 -184 -479
rect -168 -485 -165 -479
rect -156 -480 -128 -477
rect -156 -485 -152 -480
rect -193 -488 -152 -485
rect -122 -484 -119 -464
rect -52 -456 -49 -446
rect -52 -459 -26 -456
rect -122 -487 -74 -484
rect -66 -485 -63 -476
rect -44 -465 -41 -459
rect -66 -488 -43 -485
rect -35 -485 -32 -477
rect -35 -488 -26 -485
rect -99 -493 -84 -490
rect -66 -491 -63 -488
rect -35 -491 -32 -488
rect -75 -494 -63 -491
rect -75 -497 -72 -494
rect -44 -501 -41 -497
rect -85 -509 -82 -503
rect -66 -509 -63 -503
rect -54 -504 -26 -501
rect -54 -509 -50 -504
rect -91 -512 -50 -509
rect -244 -524 -202 -521
rect -339 -557 -323 -554
rect -319 -529 -293 -526
rect -416 -562 -377 -559
rect -369 -565 -366 -557
rect -339 -560 -336 -557
rect -348 -570 -345 -566
rect -358 -573 -330 -570
rect -388 -583 -385 -577
rect -358 -583 -354 -573
rect -394 -586 -354 -583
rect -394 -607 -351 -606
rect -394 -609 -330 -607
rect -388 -615 -385 -609
rect -369 -615 -366 -609
rect -354 -610 -330 -609
rect -348 -616 -345 -610
rect -379 -630 -376 -627
rect -379 -633 -366 -630
rect -394 -638 -387 -635
rect -369 -636 -366 -633
rect -369 -639 -347 -636
rect -339 -636 -336 -628
rect -319 -636 -315 -529
rect -275 -527 -272 -524
rect -244 -527 -241 -524
rect -284 -530 -272 -527
rect -284 -533 -281 -530
rect -253 -537 -250 -533
rect -294 -545 -291 -539
rect -275 -545 -272 -539
rect -263 -540 -235 -537
rect -263 -545 -259 -540
rect -300 -548 -259 -545
rect -339 -637 -315 -636
rect -339 -639 -316 -637
rect -394 -644 -377 -641
rect -369 -647 -366 -639
rect -339 -642 -336 -639
rect -348 -652 -345 -648
rect -358 -655 -330 -652
rect -388 -665 -385 -659
rect -358 -665 -354 -655
rect -394 -668 -354 -665
<< m2contact >>
rect -349 491 -342 496
rect -442 245 -434 251
rect -337 248 -332 253
rect -175 194 -170 199
rect -459 -10 -448 -1
rect -338 -96 -333 -91
rect -342 -177 -335 -171
rect -468 -356 -456 -347
rect -104 -372 -96 -363
rect -444 -474 -438 -469
rect -104 -495 -99 -490
<< metal2 >>
rect -349 319 -345 491
rect -442 315 -345 319
rect -442 251 -438 315
rect -337 199 -333 248
rect -466 195 -333 199
rect -466 -10 -459 195
rect -337 97 -333 195
rect -178 97 -175 199
rect -337 92 -174 97
rect -468 -96 -338 -91
rect -468 -347 -461 -96
rect -444 -175 -342 -171
rect -444 -469 -438 -175
rect -104 -490 -99 -372
<< m3contact >>
rect -328 126 -322 131
rect -486 -127 -477 -119
rect -333 -217 -328 -212
rect -424 -563 -416 -558
<< metal3 >>
rect -327 41 -322 126
rect -486 32 -322 41
rect -486 -119 -477 32
rect -332 -285 -328 -217
rect -424 -289 -328 -285
rect -424 -558 -420 -289
<< labels >>
rlabel metal1 -254 537 -251 540 7 c0
rlabel metal1 -316 538 -313 541 1 help_c1
rlabel metal1 -316 532 -313 535 1 g0
rlabel metal1 -354 496 -351 499 1 help_c1
rlabel metal1 -415 497 -412 500 3 carry_reg
rlabel metal1 -415 491 -412 494 3 p0
rlabel metal1 -255 522 -255 522 1 gnd!
rlabel metal1 -261 567 -261 567 5 vdd!
rlabel metal1 -295 515 -295 515 1 gnd!
rlabel metal1 -298 580 -298 580 5 vdd!
rlabel metal1 -355 481 -355 481 1 gnd!
rlabel metal1 -361 526 -361 526 5 vdd!
rlabel metal1 -391 468 -391 468 1 gnd!
rlabel metal1 -391 528 -391 528 5 vdd!
rlabel metal1 -245 157 -245 157 1 gnd!
rlabel metal1 -251 202 -251 202 5 vdd!
rlabel metal1 -285 150 -285 150 1 gnd!
rlabel metal1 -288 215 -288 215 5 vdd!
rlabel metal1 -345 116 -345 116 1 gnd!
rlabel metal1 -351 161 -351 161 5 vdd!
rlabel metal1 -381 103 -381 103 1 gnd!
rlabel metal1 -381 163 -381 163 5 vdd!
rlabel metal1 -348 238 -348 238 1 gnd!
rlabel metal1 -354 283 -354 283 5 vdd!
rlabel metal1 -384 225 -384 225 1 gnd!
rlabel metal1 -384 285 -384 285 5 vdd!
rlabel metal1 -408 248 -405 251 1 help_c1
rlabel metal1 -408 254 -405 257 1 p1
rlabel metal1 -347 253 -344 256 1 help_c21
rlabel metal1 -405 132 -402 135 1 p1
rlabel metal1 -405 126 -402 129 1 g0
rlabel metal1 -344 131 -341 134 1 help_c22
rlabel metal1 -306 167 -303 170 1 g1
rlabel metal1 -306 173 -303 176 1 help_c22
rlabel metal1 -244 172 -241 175 7 inter_c11
rlabel metal1 -245 -194 -245 -194 1 gnd!
rlabel metal1 -285 -201 -285 -201 1 gnd!
rlabel metal1 -288 -136 -288 -136 5 vdd!
rlabel metal1 -386 21 -386 21 5 vdd!
rlabel metal1 -386 -39 -386 -39 1 gnd!
rlabel metal1 -356 19 -356 19 5 vdd!
rlabel metal1 -350 -26 -350 -26 1 gnd!
rlabel metal1 -383 -101 -383 -101 5 vdd!
rlabel metal1 -383 -161 -383 -161 1 gnd!
rlabel metal1 -347 -148 -347 -148 1 gnd!
rlabel metal1 -290 -49 -290 -49 5 vdd!
rlabel metal1 -287 -114 -287 -114 1 gnd!
rlabel metal1 -253 -62 -253 -62 5 vdd!
rlabel metal1 -247 -107 -247 -107 1 gnd!
rlabel metal1 -251 -149 -251 -149 5 vdd!
rlabel metal1 -353 -103 -353 -103 5 vdd!
rlabel metal1 -346 -182 -346 -182 5 vdd!
rlabel metal1 -340 -227 -340 -227 1 gnd!
rlabel metal1 -376 -240 -376 -240 1 gnd!
rlabel metal1 -376 -180 -376 -180 5 vdd!
rlabel metal1 -144 -89 -144 -89 5 vdd!
rlabel metal1 -181 -76 -181 -76 5 vdd!
rlabel metal1 -178 -141 -178 -141 1 gnd!
rlabel metal1 -138 -134 -138 -134 1 gnd!
rlabel metal1 -410 -10 -407 -7 1 help_c21
rlabel metal1 -410 -16 -407 -13 1 p2
rlabel metal1 -349 -11 -346 -8 1 help_c31
rlabel metal1 -407 -132 -404 -129 1 help_c22
rlabel metal1 -407 -138 -404 -135 1 p2
rlabel metal1 -346 -133 -343 -130 1 help_c32
rlabel metal1 -400 -211 -397 -208 1 p2
rlabel metal1 -400 -217 -397 -214 1 g1
rlabel metal1 -339 -212 -336 -209 1 help_c33
rlabel metal1 -308 -97 -305 -94 1 g2
rlabel metal1 -246 -92 -243 -89 1 inter_c21
rlabel metal1 -244 -179 -241 -176 1 inter_c22
rlabel metal1 -199 -124 -196 -121 1 inter_c22
rlabel metal1 -199 -118 -196 -115 1 inter_c21
rlabel metal1 -137 -119 -134 -116 7 c2
rlabel metal1 -132 -479 -132 -479 1 gnd!
rlabel metal1 -172 -486 -172 -486 1 gnd!
rlabel metal1 -175 -421 -175 -421 5 vdd!
rlabel metal1 -138 -434 -138 -434 5 vdd!
rlabel metal1 -370 -525 -370 -525 5 vdd!
rlabel metal1 -370 -585 -370 -585 1 gnd!
rlabel metal1 -334 -572 -334 -572 1 gnd!
rlabel metal1 -340 -527 -340 -527 5 vdd!
rlabel metal1 -347 -448 -347 -448 5 vdd!
rlabel metal1 -245 -494 -245 -494 5 vdd!
rlabel metal1 -241 -452 -241 -452 1 gnd!
rlabel metal1 -247 -407 -247 -407 5 vdd!
rlabel metal1 -281 -459 -281 -459 1 gnd!
rlabel metal1 -284 -394 -284 -394 5 vdd!
rlabel metal1 -341 -493 -341 -493 1 gnd!
rlabel metal1 -377 -506 -377 -506 1 gnd!
rlabel metal1 -377 -446 -377 -446 5 vdd!
rlabel metal1 -344 -371 -344 -371 1 gnd!
rlabel metal1 -350 -326 -350 -326 5 vdd!
rlabel metal1 -380 -384 -380 -384 1 gnd!
rlabel metal1 -380 -324 -380 -324 5 vdd!
rlabel metal1 -282 -481 -282 -481 5 vdd!
rlabel metal1 -279 -546 -279 -546 1 gnd!
rlabel metal1 -239 -539 -239 -539 1 gnd!
rlabel metal1 -343 -356 -340 -353 1 help_c41
rlabel metal1 -404 -355 -401 -352 1 help_c31
rlabel metal1 -404 -361 -401 -358 1 p3
rlabel metal1 -401 -477 -398 -474 1 help_c32
rlabel metal1 -401 -483 -398 -480 1 p3
rlabel metal1 -340 -478 -337 -475 1 help_c42
rlabel metal1 -394 -562 -391 -559 1 help_c33
rlabel metal1 -394 -556 -391 -553 1 p3
rlabel metal1 -333 -557 -330 -554 1 help_c43
rlabel metal1 -302 -436 -299 -433 1 g3
rlabel metal1 -240 -437 -237 -434 1 inter_c31
rlabel metal1 -30 -503 -30 -503 1 gnd!
rlabel metal1 -70 -510 -70 -510 1 gnd!
rlabel metal1 -73 -445 -73 -445 5 vdd!
rlabel metal1 -36 -458 -36 -458 5 vdd!
rlabel metal1 -238 -524 -235 -521 1 inter_c32
rlabel metal1 -193 -463 -190 -460 1 inter_c31
rlabel metal1 -193 -469 -190 -466 1 inter_c32
rlabel metal1 -131 -464 -128 -461 1 inter_c33
rlabel metal1 -91 -487 -88 -484 1 inter_c33
rlabel metal1 -91 -493 -88 -490 1 help_c41
rlabel metal1 -29 -488 -26 -485 7 out_carry
rlabel metal1 -137 244 -137 244 5 vdd!
rlabel metal1 -134 179 -134 179 1 gnd!
rlabel metal1 -100 231 -100 231 5 vdd!
rlabel metal1 -94 186 -94 186 1 gnd!
rlabel metal1 -155 202 -152 205 1 inter_c11
rlabel metal1 -93 201 -90 204 7 c1
rlabel metal1 -155 196 -152 199 1 help_c21
rlabel metal1 -308 -91 -305 -88 1 help_c31
rlabel metal1 -306 -178 -303 -175 1 help_c32
rlabel metal1 -306 -184 -303 -181 1 help_c33
rlabel metal1 -370 -607 -370 -607 5 vdd!
rlabel metal1 -370 -667 -370 -667 1 gnd!
rlabel metal1 -334 -654 -334 -654 1 gnd!
rlabel metal1 -340 -609 -340 -609 5 vdd!
rlabel metal1 -394 -644 -391 -641 1 g2
rlabel metal1 -394 -638 -391 -635 1 p3
rlabel metal1 -333 -639 -330 -636 1 help_c44
rlabel metal1 -302 -442 -299 -439 1 help_c42
rlabel metal1 -300 -523 -297 -520 1 help_c43
rlabel metal1 -300 -529 -297 -526 1 help_c44
<< end >>
